magic
tech sky130B
magscale 1 2
timestamp 1659562972
<< obsli1 >>
rect 1104 2159 278852 357425
<< obsm1 >>
rect 14 2128 279666 357456
<< metal2 >>
rect 18 359200 74 360000
rect 662 359200 718 360000
rect 1306 359200 1362 360000
rect 1950 359200 2006 360000
rect 2594 359200 2650 360000
rect 3238 359200 3294 360000
rect 3882 359200 3938 360000
rect 4526 359200 4582 360000
rect 5170 359200 5226 360000
rect 6458 359200 6514 360000
rect 7102 359200 7158 360000
rect 7746 359200 7802 360000
rect 8390 359200 8446 360000
rect 9034 359200 9090 360000
rect 9678 359200 9734 360000
rect 10322 359200 10378 360000
rect 10966 359200 11022 360000
rect 12254 359200 12310 360000
rect 12898 359200 12954 360000
rect 13542 359200 13598 360000
rect 14186 359200 14242 360000
rect 14830 359200 14886 360000
rect 15474 359200 15530 360000
rect 16118 359200 16174 360000
rect 16762 359200 16818 360000
rect 17406 359200 17462 360000
rect 18694 359200 18750 360000
rect 19338 359200 19394 360000
rect 19982 359200 20038 360000
rect 20626 359200 20682 360000
rect 21270 359200 21326 360000
rect 21914 359200 21970 360000
rect 22558 359200 22614 360000
rect 23202 359200 23258 360000
rect 24490 359200 24546 360000
rect 25134 359200 25190 360000
rect 25778 359200 25834 360000
rect 26422 359200 26478 360000
rect 27066 359200 27122 360000
rect 27710 359200 27766 360000
rect 28354 359200 28410 360000
rect 28998 359200 29054 360000
rect 29642 359200 29698 360000
rect 30930 359200 30986 360000
rect 31574 359200 31630 360000
rect 32218 359200 32274 360000
rect 32862 359200 32918 360000
rect 33506 359200 33562 360000
rect 34150 359200 34206 360000
rect 34794 359200 34850 360000
rect 35438 359200 35494 360000
rect 36726 359200 36782 360000
rect 37370 359200 37426 360000
rect 38014 359200 38070 360000
rect 38658 359200 38714 360000
rect 39302 359200 39358 360000
rect 39946 359200 40002 360000
rect 40590 359200 40646 360000
rect 41234 359200 41290 360000
rect 41878 359200 41934 360000
rect 43166 359200 43222 360000
rect 43810 359200 43866 360000
rect 44454 359200 44510 360000
rect 45098 359200 45154 360000
rect 45742 359200 45798 360000
rect 46386 359200 46442 360000
rect 47030 359200 47086 360000
rect 47674 359200 47730 360000
rect 48962 359200 49018 360000
rect 49606 359200 49662 360000
rect 50250 359200 50306 360000
rect 50894 359200 50950 360000
rect 51538 359200 51594 360000
rect 52182 359200 52238 360000
rect 52826 359200 52882 360000
rect 53470 359200 53526 360000
rect 54758 359200 54814 360000
rect 55402 359200 55458 360000
rect 56046 359200 56102 360000
rect 56690 359200 56746 360000
rect 57334 359200 57390 360000
rect 57978 359200 58034 360000
rect 58622 359200 58678 360000
rect 59266 359200 59322 360000
rect 59910 359200 59966 360000
rect 61198 359200 61254 360000
rect 61842 359200 61898 360000
rect 62486 359200 62542 360000
rect 63130 359200 63186 360000
rect 63774 359200 63830 360000
rect 64418 359200 64474 360000
rect 65062 359200 65118 360000
rect 65706 359200 65762 360000
rect 66994 359200 67050 360000
rect 67638 359200 67694 360000
rect 68282 359200 68338 360000
rect 68926 359200 68982 360000
rect 69570 359200 69626 360000
rect 70214 359200 70270 360000
rect 70858 359200 70914 360000
rect 71502 359200 71558 360000
rect 72146 359200 72202 360000
rect 73434 359200 73490 360000
rect 74078 359200 74134 360000
rect 74722 359200 74778 360000
rect 75366 359200 75422 360000
rect 76010 359200 76066 360000
rect 76654 359200 76710 360000
rect 77298 359200 77354 360000
rect 77942 359200 77998 360000
rect 79230 359200 79286 360000
rect 79874 359200 79930 360000
rect 80518 359200 80574 360000
rect 81162 359200 81218 360000
rect 81806 359200 81862 360000
rect 82450 359200 82506 360000
rect 83094 359200 83150 360000
rect 83738 359200 83794 360000
rect 84382 359200 84438 360000
rect 85670 359200 85726 360000
rect 86314 359200 86370 360000
rect 86958 359200 87014 360000
rect 87602 359200 87658 360000
rect 88246 359200 88302 360000
rect 88890 359200 88946 360000
rect 89534 359200 89590 360000
rect 90178 359200 90234 360000
rect 91466 359200 91522 360000
rect 92110 359200 92166 360000
rect 92754 359200 92810 360000
rect 93398 359200 93454 360000
rect 94042 359200 94098 360000
rect 94686 359200 94742 360000
rect 95330 359200 95386 360000
rect 95974 359200 96030 360000
rect 96618 359200 96674 360000
rect 97906 359200 97962 360000
rect 98550 359200 98606 360000
rect 99194 359200 99250 360000
rect 99838 359200 99894 360000
rect 100482 359200 100538 360000
rect 101126 359200 101182 360000
rect 101770 359200 101826 360000
rect 102414 359200 102470 360000
rect 103702 359200 103758 360000
rect 104346 359200 104402 360000
rect 104990 359200 105046 360000
rect 105634 359200 105690 360000
rect 106278 359200 106334 360000
rect 106922 359200 106978 360000
rect 107566 359200 107622 360000
rect 108210 359200 108266 360000
rect 108854 359200 108910 360000
rect 110142 359200 110198 360000
rect 110786 359200 110842 360000
rect 111430 359200 111486 360000
rect 112074 359200 112130 360000
rect 112718 359200 112774 360000
rect 113362 359200 113418 360000
rect 114006 359200 114062 360000
rect 114650 359200 114706 360000
rect 115938 359200 115994 360000
rect 116582 359200 116638 360000
rect 117226 359200 117282 360000
rect 117870 359200 117926 360000
rect 118514 359200 118570 360000
rect 119158 359200 119214 360000
rect 119802 359200 119858 360000
rect 120446 359200 120502 360000
rect 121090 359200 121146 360000
rect 122378 359200 122434 360000
rect 123022 359200 123078 360000
rect 123666 359200 123722 360000
rect 124310 359200 124366 360000
rect 124954 359200 125010 360000
rect 125598 359200 125654 360000
rect 126242 359200 126298 360000
rect 126886 359200 126942 360000
rect 128174 359200 128230 360000
rect 128818 359200 128874 360000
rect 129462 359200 129518 360000
rect 130106 359200 130162 360000
rect 130750 359200 130806 360000
rect 131394 359200 131450 360000
rect 132038 359200 132094 360000
rect 132682 359200 132738 360000
rect 133970 359200 134026 360000
rect 134614 359200 134670 360000
rect 135258 359200 135314 360000
rect 135902 359200 135958 360000
rect 136546 359200 136602 360000
rect 137190 359200 137246 360000
rect 137834 359200 137890 360000
rect 138478 359200 138534 360000
rect 139122 359200 139178 360000
rect 140410 359200 140466 360000
rect 141054 359200 141110 360000
rect 141698 359200 141754 360000
rect 142342 359200 142398 360000
rect 142986 359200 143042 360000
rect 143630 359200 143686 360000
rect 144274 359200 144330 360000
rect 144918 359200 144974 360000
rect 146206 359200 146262 360000
rect 146850 359200 146906 360000
rect 147494 359200 147550 360000
rect 148138 359200 148194 360000
rect 148782 359200 148838 360000
rect 149426 359200 149482 360000
rect 150070 359200 150126 360000
rect 150714 359200 150770 360000
rect 151358 359200 151414 360000
rect 152646 359200 152702 360000
rect 153290 359200 153346 360000
rect 153934 359200 153990 360000
rect 154578 359200 154634 360000
rect 155222 359200 155278 360000
rect 155866 359200 155922 360000
rect 156510 359200 156566 360000
rect 157154 359200 157210 360000
rect 158442 359200 158498 360000
rect 159086 359200 159142 360000
rect 159730 359200 159786 360000
rect 160374 359200 160430 360000
rect 161018 359200 161074 360000
rect 161662 359200 161718 360000
rect 162306 359200 162362 360000
rect 162950 359200 163006 360000
rect 163594 359200 163650 360000
rect 164882 359200 164938 360000
rect 165526 359200 165582 360000
rect 166170 359200 166226 360000
rect 166814 359200 166870 360000
rect 167458 359200 167514 360000
rect 168102 359200 168158 360000
rect 168746 359200 168802 360000
rect 169390 359200 169446 360000
rect 170678 359200 170734 360000
rect 171322 359200 171378 360000
rect 171966 359200 172022 360000
rect 172610 359200 172666 360000
rect 173254 359200 173310 360000
rect 173898 359200 173954 360000
rect 174542 359200 174598 360000
rect 175186 359200 175242 360000
rect 175830 359200 175886 360000
rect 177118 359200 177174 360000
rect 177762 359200 177818 360000
rect 178406 359200 178462 360000
rect 179050 359200 179106 360000
rect 179694 359200 179750 360000
rect 180338 359200 180394 360000
rect 180982 359200 181038 360000
rect 181626 359200 181682 360000
rect 182914 359200 182970 360000
rect 183558 359200 183614 360000
rect 184202 359200 184258 360000
rect 184846 359200 184902 360000
rect 185490 359200 185546 360000
rect 186134 359200 186190 360000
rect 186778 359200 186834 360000
rect 187422 359200 187478 360000
rect 188066 359200 188122 360000
rect 189354 359200 189410 360000
rect 189998 359200 190054 360000
rect 190642 359200 190698 360000
rect 191286 359200 191342 360000
rect 191930 359200 191986 360000
rect 192574 359200 192630 360000
rect 193218 359200 193274 360000
rect 193862 359200 193918 360000
rect 195150 359200 195206 360000
rect 195794 359200 195850 360000
rect 196438 359200 196494 360000
rect 197082 359200 197138 360000
rect 197726 359200 197782 360000
rect 198370 359200 198426 360000
rect 199014 359200 199070 360000
rect 199658 359200 199714 360000
rect 200302 359200 200358 360000
rect 201590 359200 201646 360000
rect 202234 359200 202290 360000
rect 202878 359200 202934 360000
rect 203522 359200 203578 360000
rect 204166 359200 204222 360000
rect 204810 359200 204866 360000
rect 205454 359200 205510 360000
rect 206098 359200 206154 360000
rect 207386 359200 207442 360000
rect 208030 359200 208086 360000
rect 208674 359200 208730 360000
rect 209318 359200 209374 360000
rect 209962 359200 210018 360000
rect 210606 359200 210662 360000
rect 211250 359200 211306 360000
rect 211894 359200 211950 360000
rect 213182 359200 213238 360000
rect 213826 359200 213882 360000
rect 214470 359200 214526 360000
rect 215114 359200 215170 360000
rect 215758 359200 215814 360000
rect 216402 359200 216458 360000
rect 217046 359200 217102 360000
rect 217690 359200 217746 360000
rect 218334 359200 218390 360000
rect 219622 359200 219678 360000
rect 220266 359200 220322 360000
rect 220910 359200 220966 360000
rect 221554 359200 221610 360000
rect 222198 359200 222254 360000
rect 222842 359200 222898 360000
rect 223486 359200 223542 360000
rect 224130 359200 224186 360000
rect 225418 359200 225474 360000
rect 226062 359200 226118 360000
rect 226706 359200 226762 360000
rect 227350 359200 227406 360000
rect 227994 359200 228050 360000
rect 228638 359200 228694 360000
rect 229282 359200 229338 360000
rect 229926 359200 229982 360000
rect 230570 359200 230626 360000
rect 231858 359200 231914 360000
rect 232502 359200 232558 360000
rect 233146 359200 233202 360000
rect 233790 359200 233846 360000
rect 234434 359200 234490 360000
rect 235078 359200 235134 360000
rect 235722 359200 235778 360000
rect 236366 359200 236422 360000
rect 237654 359200 237710 360000
rect 238298 359200 238354 360000
rect 238942 359200 238998 360000
rect 239586 359200 239642 360000
rect 240230 359200 240286 360000
rect 240874 359200 240930 360000
rect 241518 359200 241574 360000
rect 242162 359200 242218 360000
rect 242806 359200 242862 360000
rect 244094 359200 244150 360000
rect 244738 359200 244794 360000
rect 245382 359200 245438 360000
rect 246026 359200 246082 360000
rect 246670 359200 246726 360000
rect 247314 359200 247370 360000
rect 247958 359200 248014 360000
rect 248602 359200 248658 360000
rect 249890 359200 249946 360000
rect 250534 359200 250590 360000
rect 251178 359200 251234 360000
rect 251822 359200 251878 360000
rect 252466 359200 252522 360000
rect 253110 359200 253166 360000
rect 253754 359200 253810 360000
rect 254398 359200 254454 360000
rect 255042 359200 255098 360000
rect 256330 359200 256386 360000
rect 256974 359200 257030 360000
rect 257618 359200 257674 360000
rect 258262 359200 258318 360000
rect 258906 359200 258962 360000
rect 259550 359200 259606 360000
rect 260194 359200 260250 360000
rect 260838 359200 260894 360000
rect 262126 359200 262182 360000
rect 262770 359200 262826 360000
rect 263414 359200 263470 360000
rect 264058 359200 264114 360000
rect 264702 359200 264758 360000
rect 265346 359200 265402 360000
rect 265990 359200 266046 360000
rect 266634 359200 266690 360000
rect 267278 359200 267334 360000
rect 268566 359200 268622 360000
rect 269210 359200 269266 360000
rect 269854 359200 269910 360000
rect 270498 359200 270554 360000
rect 271142 359200 271198 360000
rect 271786 359200 271842 360000
rect 272430 359200 272486 360000
rect 273074 359200 273130 360000
rect 274362 359200 274418 360000
rect 275006 359200 275062 360000
rect 275650 359200 275706 360000
rect 276294 359200 276350 360000
rect 276938 359200 276994 360000
rect 277582 359200 277638 360000
rect 278226 359200 278282 360000
rect 278870 359200 278926 360000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 48962 0 49018 800
rect 49606 0 49662 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 53470 0 53526 800
rect 54114 0 54170 800
rect 55402 0 55458 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59266 0 59322 800
rect 59910 0 59966 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65062 0 65118 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74722 0 74778 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 76654 0 76710 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80518 0 80574 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82450 0 82506 800
rect 83094 0 83150 800
rect 83738 0 83794 800
rect 84382 0 84438 800
rect 85670 0 85726 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 87602 0 87658 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 89534 0 89590 800
rect 90178 0 90234 800
rect 91466 0 91522 800
rect 92110 0 92166 800
rect 92754 0 92810 800
rect 93398 0 93454 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95330 0 95386 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99194 0 99250 800
rect 99838 0 99894 800
rect 100482 0 100538 800
rect 101126 0 101182 800
rect 101770 0 101826 800
rect 102414 0 102470 800
rect 103702 0 103758 800
rect 104346 0 104402 800
rect 104990 0 105046 800
rect 105634 0 105690 800
rect 106278 0 106334 800
rect 106922 0 106978 800
rect 107566 0 107622 800
rect 108210 0 108266 800
rect 108854 0 108910 800
rect 110142 0 110198 800
rect 110786 0 110842 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 112718 0 112774 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 114650 0 114706 800
rect 115938 0 115994 800
rect 116582 0 116638 800
rect 117226 0 117282 800
rect 117870 0 117926 800
rect 118514 0 118570 800
rect 119158 0 119214 800
rect 119802 0 119858 800
rect 120446 0 120502 800
rect 121090 0 121146 800
rect 122378 0 122434 800
rect 123022 0 123078 800
rect 123666 0 123722 800
rect 124310 0 124366 800
rect 124954 0 125010 800
rect 125598 0 125654 800
rect 126242 0 126298 800
rect 126886 0 126942 800
rect 128174 0 128230 800
rect 128818 0 128874 800
rect 129462 0 129518 800
rect 130106 0 130162 800
rect 130750 0 130806 800
rect 131394 0 131450 800
rect 132038 0 132094 800
rect 132682 0 132738 800
rect 133326 0 133382 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 135902 0 135958 800
rect 136546 0 136602 800
rect 137190 0 137246 800
rect 137834 0 137890 800
rect 138478 0 138534 800
rect 139122 0 139178 800
rect 140410 0 140466 800
rect 141054 0 141110 800
rect 141698 0 141754 800
rect 142342 0 142398 800
rect 142986 0 143042 800
rect 143630 0 143686 800
rect 144274 0 144330 800
rect 144918 0 144974 800
rect 145562 0 145618 800
rect 146850 0 146906 800
rect 147494 0 147550 800
rect 148138 0 148194 800
rect 148782 0 148838 800
rect 149426 0 149482 800
rect 150070 0 150126 800
rect 150714 0 150770 800
rect 151358 0 151414 800
rect 152646 0 152702 800
rect 153290 0 153346 800
rect 153934 0 153990 800
rect 154578 0 154634 800
rect 155222 0 155278 800
rect 155866 0 155922 800
rect 156510 0 156566 800
rect 157154 0 157210 800
rect 158442 0 158498 800
rect 159086 0 159142 800
rect 159730 0 159786 800
rect 160374 0 160430 800
rect 161018 0 161074 800
rect 161662 0 161718 800
rect 162306 0 162362 800
rect 162950 0 163006 800
rect 163594 0 163650 800
rect 164882 0 164938 800
rect 165526 0 165582 800
rect 166170 0 166226 800
rect 166814 0 166870 800
rect 167458 0 167514 800
rect 168102 0 168158 800
rect 168746 0 168802 800
rect 169390 0 169446 800
rect 170678 0 170734 800
rect 171322 0 171378 800
rect 171966 0 172022 800
rect 172610 0 172666 800
rect 173254 0 173310 800
rect 173898 0 173954 800
rect 174542 0 174598 800
rect 175186 0 175242 800
rect 175830 0 175886 800
rect 177118 0 177174 800
rect 177762 0 177818 800
rect 178406 0 178462 800
rect 179050 0 179106 800
rect 179694 0 179750 800
rect 180338 0 180394 800
rect 180982 0 181038 800
rect 181626 0 181682 800
rect 182914 0 182970 800
rect 183558 0 183614 800
rect 184202 0 184258 800
rect 184846 0 184902 800
rect 185490 0 185546 800
rect 186134 0 186190 800
rect 186778 0 186834 800
rect 187422 0 187478 800
rect 188066 0 188122 800
rect 189354 0 189410 800
rect 189998 0 190054 800
rect 190642 0 190698 800
rect 191286 0 191342 800
rect 191930 0 191986 800
rect 192574 0 192630 800
rect 193218 0 193274 800
rect 193862 0 193918 800
rect 195150 0 195206 800
rect 195794 0 195850 800
rect 196438 0 196494 800
rect 197082 0 197138 800
rect 197726 0 197782 800
rect 198370 0 198426 800
rect 199014 0 199070 800
rect 199658 0 199714 800
rect 200302 0 200358 800
rect 201590 0 201646 800
rect 202234 0 202290 800
rect 202878 0 202934 800
rect 203522 0 203578 800
rect 204166 0 204222 800
rect 204810 0 204866 800
rect 205454 0 205510 800
rect 206098 0 206154 800
rect 207386 0 207442 800
rect 208030 0 208086 800
rect 208674 0 208730 800
rect 209318 0 209374 800
rect 209962 0 210018 800
rect 210606 0 210662 800
rect 211250 0 211306 800
rect 211894 0 211950 800
rect 212538 0 212594 800
rect 213826 0 213882 800
rect 214470 0 214526 800
rect 215114 0 215170 800
rect 215758 0 215814 800
rect 216402 0 216458 800
rect 217046 0 217102 800
rect 217690 0 217746 800
rect 218334 0 218390 800
rect 219622 0 219678 800
rect 220266 0 220322 800
rect 220910 0 220966 800
rect 221554 0 221610 800
rect 222198 0 222254 800
rect 222842 0 222898 800
rect 223486 0 223542 800
rect 224130 0 224186 800
rect 224774 0 224830 800
rect 226062 0 226118 800
rect 226706 0 226762 800
rect 227350 0 227406 800
rect 227994 0 228050 800
rect 228638 0 228694 800
rect 229282 0 229338 800
rect 229926 0 229982 800
rect 230570 0 230626 800
rect 231858 0 231914 800
rect 232502 0 232558 800
rect 233146 0 233202 800
rect 233790 0 233846 800
rect 234434 0 234490 800
rect 235078 0 235134 800
rect 235722 0 235778 800
rect 236366 0 236422 800
rect 237654 0 237710 800
rect 238298 0 238354 800
rect 238942 0 238998 800
rect 239586 0 239642 800
rect 240230 0 240286 800
rect 240874 0 240930 800
rect 241518 0 241574 800
rect 242162 0 242218 800
rect 242806 0 242862 800
rect 244094 0 244150 800
rect 244738 0 244794 800
rect 245382 0 245438 800
rect 246026 0 246082 800
rect 246670 0 246726 800
rect 247314 0 247370 800
rect 247958 0 248014 800
rect 248602 0 248658 800
rect 249890 0 249946 800
rect 250534 0 250590 800
rect 251178 0 251234 800
rect 251822 0 251878 800
rect 252466 0 252522 800
rect 253110 0 253166 800
rect 253754 0 253810 800
rect 254398 0 254454 800
rect 255042 0 255098 800
rect 256330 0 256386 800
rect 256974 0 257030 800
rect 257618 0 257674 800
rect 258262 0 258318 800
rect 258906 0 258962 800
rect 259550 0 259606 800
rect 260194 0 260250 800
rect 260838 0 260894 800
rect 262126 0 262182 800
rect 262770 0 262826 800
rect 263414 0 263470 800
rect 264058 0 264114 800
rect 264702 0 264758 800
rect 265346 0 265402 800
rect 265990 0 266046 800
rect 266634 0 266690 800
rect 267278 0 267334 800
rect 268566 0 268622 800
rect 269210 0 269266 800
rect 269854 0 269910 800
rect 270498 0 270554 800
rect 271142 0 271198 800
rect 271786 0 271842 800
rect 272430 0 272486 800
rect 273074 0 273130 800
rect 274362 0 274418 800
rect 275006 0 275062 800
rect 275650 0 275706 800
rect 276294 0 276350 800
rect 276938 0 276994 800
rect 277582 0 277638 800
rect 278226 0 278282 800
rect 278870 0 278926 800
rect 279514 0 279570 800
<< obsm2 >>
rect 130 359144 606 359258
rect 774 359144 1250 359258
rect 1418 359144 1894 359258
rect 2062 359144 2538 359258
rect 2706 359144 3182 359258
rect 3350 359144 3826 359258
rect 3994 359144 4470 359258
rect 4638 359144 5114 359258
rect 5282 359144 6402 359258
rect 6570 359144 7046 359258
rect 7214 359144 7690 359258
rect 7858 359144 8334 359258
rect 8502 359144 8978 359258
rect 9146 359144 9622 359258
rect 9790 359144 10266 359258
rect 10434 359144 10910 359258
rect 11078 359144 12198 359258
rect 12366 359144 12842 359258
rect 13010 359144 13486 359258
rect 13654 359144 14130 359258
rect 14298 359144 14774 359258
rect 14942 359144 15418 359258
rect 15586 359144 16062 359258
rect 16230 359144 16706 359258
rect 16874 359144 17350 359258
rect 17518 359144 18638 359258
rect 18806 359144 19282 359258
rect 19450 359144 19926 359258
rect 20094 359144 20570 359258
rect 20738 359144 21214 359258
rect 21382 359144 21858 359258
rect 22026 359144 22502 359258
rect 22670 359144 23146 359258
rect 23314 359144 24434 359258
rect 24602 359144 25078 359258
rect 25246 359144 25722 359258
rect 25890 359144 26366 359258
rect 26534 359144 27010 359258
rect 27178 359144 27654 359258
rect 27822 359144 28298 359258
rect 28466 359144 28942 359258
rect 29110 359144 29586 359258
rect 29754 359144 30874 359258
rect 31042 359144 31518 359258
rect 31686 359144 32162 359258
rect 32330 359144 32806 359258
rect 32974 359144 33450 359258
rect 33618 359144 34094 359258
rect 34262 359144 34738 359258
rect 34906 359144 35382 359258
rect 35550 359144 36670 359258
rect 36838 359144 37314 359258
rect 37482 359144 37958 359258
rect 38126 359144 38602 359258
rect 38770 359144 39246 359258
rect 39414 359144 39890 359258
rect 40058 359144 40534 359258
rect 40702 359144 41178 359258
rect 41346 359144 41822 359258
rect 41990 359144 43110 359258
rect 43278 359144 43754 359258
rect 43922 359144 44398 359258
rect 44566 359144 45042 359258
rect 45210 359144 45686 359258
rect 45854 359144 46330 359258
rect 46498 359144 46974 359258
rect 47142 359144 47618 359258
rect 47786 359144 48906 359258
rect 49074 359144 49550 359258
rect 49718 359144 50194 359258
rect 50362 359144 50838 359258
rect 51006 359144 51482 359258
rect 51650 359144 52126 359258
rect 52294 359144 52770 359258
rect 52938 359144 53414 359258
rect 53582 359144 54702 359258
rect 54870 359144 55346 359258
rect 55514 359144 55990 359258
rect 56158 359144 56634 359258
rect 56802 359144 57278 359258
rect 57446 359144 57922 359258
rect 58090 359144 58566 359258
rect 58734 359144 59210 359258
rect 59378 359144 59854 359258
rect 60022 359144 61142 359258
rect 61310 359144 61786 359258
rect 61954 359144 62430 359258
rect 62598 359144 63074 359258
rect 63242 359144 63718 359258
rect 63886 359144 64362 359258
rect 64530 359144 65006 359258
rect 65174 359144 65650 359258
rect 65818 359144 66938 359258
rect 67106 359144 67582 359258
rect 67750 359144 68226 359258
rect 68394 359144 68870 359258
rect 69038 359144 69514 359258
rect 69682 359144 70158 359258
rect 70326 359144 70802 359258
rect 70970 359144 71446 359258
rect 71614 359144 72090 359258
rect 72258 359144 73378 359258
rect 73546 359144 74022 359258
rect 74190 359144 74666 359258
rect 74834 359144 75310 359258
rect 75478 359144 75954 359258
rect 76122 359144 76598 359258
rect 76766 359144 77242 359258
rect 77410 359144 77886 359258
rect 78054 359144 79174 359258
rect 79342 359144 79818 359258
rect 79986 359144 80462 359258
rect 80630 359144 81106 359258
rect 81274 359144 81750 359258
rect 81918 359144 82394 359258
rect 82562 359144 83038 359258
rect 83206 359144 83682 359258
rect 83850 359144 84326 359258
rect 84494 359144 85614 359258
rect 85782 359144 86258 359258
rect 86426 359144 86902 359258
rect 87070 359144 87546 359258
rect 87714 359144 88190 359258
rect 88358 359144 88834 359258
rect 89002 359144 89478 359258
rect 89646 359144 90122 359258
rect 90290 359144 91410 359258
rect 91578 359144 92054 359258
rect 92222 359144 92698 359258
rect 92866 359144 93342 359258
rect 93510 359144 93986 359258
rect 94154 359144 94630 359258
rect 94798 359144 95274 359258
rect 95442 359144 95918 359258
rect 96086 359144 96562 359258
rect 96730 359144 97850 359258
rect 98018 359144 98494 359258
rect 98662 359144 99138 359258
rect 99306 359144 99782 359258
rect 99950 359144 100426 359258
rect 100594 359144 101070 359258
rect 101238 359144 101714 359258
rect 101882 359144 102358 359258
rect 102526 359144 103646 359258
rect 103814 359144 104290 359258
rect 104458 359144 104934 359258
rect 105102 359144 105578 359258
rect 105746 359144 106222 359258
rect 106390 359144 106866 359258
rect 107034 359144 107510 359258
rect 107678 359144 108154 359258
rect 108322 359144 108798 359258
rect 108966 359144 110086 359258
rect 110254 359144 110730 359258
rect 110898 359144 111374 359258
rect 111542 359144 112018 359258
rect 112186 359144 112662 359258
rect 112830 359144 113306 359258
rect 113474 359144 113950 359258
rect 114118 359144 114594 359258
rect 114762 359144 115882 359258
rect 116050 359144 116526 359258
rect 116694 359144 117170 359258
rect 117338 359144 117814 359258
rect 117982 359144 118458 359258
rect 118626 359144 119102 359258
rect 119270 359144 119746 359258
rect 119914 359144 120390 359258
rect 120558 359144 121034 359258
rect 121202 359144 122322 359258
rect 122490 359144 122966 359258
rect 123134 359144 123610 359258
rect 123778 359144 124254 359258
rect 124422 359144 124898 359258
rect 125066 359144 125542 359258
rect 125710 359144 126186 359258
rect 126354 359144 126830 359258
rect 126998 359144 128118 359258
rect 128286 359144 128762 359258
rect 128930 359144 129406 359258
rect 129574 359144 130050 359258
rect 130218 359144 130694 359258
rect 130862 359144 131338 359258
rect 131506 359144 131982 359258
rect 132150 359144 132626 359258
rect 132794 359144 133914 359258
rect 134082 359144 134558 359258
rect 134726 359144 135202 359258
rect 135370 359144 135846 359258
rect 136014 359144 136490 359258
rect 136658 359144 137134 359258
rect 137302 359144 137778 359258
rect 137946 359144 138422 359258
rect 138590 359144 139066 359258
rect 139234 359144 140354 359258
rect 140522 359144 140998 359258
rect 141166 359144 141642 359258
rect 141810 359144 142286 359258
rect 142454 359144 142930 359258
rect 143098 359144 143574 359258
rect 143742 359144 144218 359258
rect 144386 359144 144862 359258
rect 145030 359144 146150 359258
rect 146318 359144 146794 359258
rect 146962 359144 147438 359258
rect 147606 359144 148082 359258
rect 148250 359144 148726 359258
rect 148894 359144 149370 359258
rect 149538 359144 150014 359258
rect 150182 359144 150658 359258
rect 150826 359144 151302 359258
rect 151470 359144 152590 359258
rect 152758 359144 153234 359258
rect 153402 359144 153878 359258
rect 154046 359144 154522 359258
rect 154690 359144 155166 359258
rect 155334 359144 155810 359258
rect 155978 359144 156454 359258
rect 156622 359144 157098 359258
rect 157266 359144 158386 359258
rect 158554 359144 159030 359258
rect 159198 359144 159674 359258
rect 159842 359144 160318 359258
rect 160486 359144 160962 359258
rect 161130 359144 161606 359258
rect 161774 359144 162250 359258
rect 162418 359144 162894 359258
rect 163062 359144 163538 359258
rect 163706 359144 164826 359258
rect 164994 359144 165470 359258
rect 165638 359144 166114 359258
rect 166282 359144 166758 359258
rect 166926 359144 167402 359258
rect 167570 359144 168046 359258
rect 168214 359144 168690 359258
rect 168858 359144 169334 359258
rect 169502 359144 170622 359258
rect 170790 359144 171266 359258
rect 171434 359144 171910 359258
rect 172078 359144 172554 359258
rect 172722 359144 173198 359258
rect 173366 359144 173842 359258
rect 174010 359144 174486 359258
rect 174654 359144 175130 359258
rect 175298 359144 175774 359258
rect 175942 359144 177062 359258
rect 177230 359144 177706 359258
rect 177874 359144 178350 359258
rect 178518 359144 178994 359258
rect 179162 359144 179638 359258
rect 179806 359144 180282 359258
rect 180450 359144 180926 359258
rect 181094 359144 181570 359258
rect 181738 359144 182858 359258
rect 183026 359144 183502 359258
rect 183670 359144 184146 359258
rect 184314 359144 184790 359258
rect 184958 359144 185434 359258
rect 185602 359144 186078 359258
rect 186246 359144 186722 359258
rect 186890 359144 187366 359258
rect 187534 359144 188010 359258
rect 188178 359144 189298 359258
rect 189466 359144 189942 359258
rect 190110 359144 190586 359258
rect 190754 359144 191230 359258
rect 191398 359144 191874 359258
rect 192042 359144 192518 359258
rect 192686 359144 193162 359258
rect 193330 359144 193806 359258
rect 193974 359144 195094 359258
rect 195262 359144 195738 359258
rect 195906 359144 196382 359258
rect 196550 359144 197026 359258
rect 197194 359144 197670 359258
rect 197838 359144 198314 359258
rect 198482 359144 198958 359258
rect 199126 359144 199602 359258
rect 199770 359144 200246 359258
rect 200414 359144 201534 359258
rect 201702 359144 202178 359258
rect 202346 359144 202822 359258
rect 202990 359144 203466 359258
rect 203634 359144 204110 359258
rect 204278 359144 204754 359258
rect 204922 359144 205398 359258
rect 205566 359144 206042 359258
rect 206210 359144 207330 359258
rect 207498 359144 207974 359258
rect 208142 359144 208618 359258
rect 208786 359144 209262 359258
rect 209430 359144 209906 359258
rect 210074 359144 210550 359258
rect 210718 359144 211194 359258
rect 211362 359144 211838 359258
rect 212006 359144 213126 359258
rect 213294 359144 213770 359258
rect 213938 359144 214414 359258
rect 214582 359144 215058 359258
rect 215226 359144 215702 359258
rect 215870 359144 216346 359258
rect 216514 359144 216990 359258
rect 217158 359144 217634 359258
rect 217802 359144 218278 359258
rect 218446 359144 219566 359258
rect 219734 359144 220210 359258
rect 220378 359144 220854 359258
rect 221022 359144 221498 359258
rect 221666 359144 222142 359258
rect 222310 359144 222786 359258
rect 222954 359144 223430 359258
rect 223598 359144 224074 359258
rect 224242 359144 225362 359258
rect 225530 359144 226006 359258
rect 226174 359144 226650 359258
rect 226818 359144 227294 359258
rect 227462 359144 227938 359258
rect 228106 359144 228582 359258
rect 228750 359144 229226 359258
rect 229394 359144 229870 359258
rect 230038 359144 230514 359258
rect 230682 359144 231802 359258
rect 231970 359144 232446 359258
rect 232614 359144 233090 359258
rect 233258 359144 233734 359258
rect 233902 359144 234378 359258
rect 234546 359144 235022 359258
rect 235190 359144 235666 359258
rect 235834 359144 236310 359258
rect 236478 359144 237598 359258
rect 237766 359144 238242 359258
rect 238410 359144 238886 359258
rect 239054 359144 239530 359258
rect 239698 359144 240174 359258
rect 240342 359144 240818 359258
rect 240986 359144 241462 359258
rect 241630 359144 242106 359258
rect 242274 359144 242750 359258
rect 242918 359144 244038 359258
rect 244206 359144 244682 359258
rect 244850 359144 245326 359258
rect 245494 359144 245970 359258
rect 246138 359144 246614 359258
rect 246782 359144 247258 359258
rect 247426 359144 247902 359258
rect 248070 359144 248546 359258
rect 248714 359144 249834 359258
rect 250002 359144 250478 359258
rect 250646 359144 251122 359258
rect 251290 359144 251766 359258
rect 251934 359144 252410 359258
rect 252578 359144 253054 359258
rect 253222 359144 253698 359258
rect 253866 359144 254342 359258
rect 254510 359144 254986 359258
rect 255154 359144 256274 359258
rect 256442 359144 256918 359258
rect 257086 359144 257562 359258
rect 257730 359144 258206 359258
rect 258374 359144 258850 359258
rect 259018 359144 259494 359258
rect 259662 359144 260138 359258
rect 260306 359144 260782 359258
rect 260950 359144 262070 359258
rect 262238 359144 262714 359258
rect 262882 359144 263358 359258
rect 263526 359144 264002 359258
rect 264170 359144 264646 359258
rect 264814 359144 265290 359258
rect 265458 359144 265934 359258
rect 266102 359144 266578 359258
rect 266746 359144 267222 359258
rect 267390 359144 268510 359258
rect 268678 359144 269154 359258
rect 269322 359144 269798 359258
rect 269966 359144 270442 359258
rect 270610 359144 271086 359258
rect 271254 359144 271730 359258
rect 271898 359144 272374 359258
rect 272542 359144 273018 359258
rect 273186 359144 274306 359258
rect 274474 359144 274950 359258
rect 275118 359144 275594 359258
rect 275762 359144 276238 359258
rect 276406 359144 276882 359258
rect 277050 359144 277526 359258
rect 277694 359144 278170 359258
rect 278338 359144 278814 359258
rect 278982 359144 279660 359258
rect 20 856 279660 359144
rect 130 711 606 856
rect 774 711 1250 856
rect 1418 711 1894 856
rect 2062 711 2538 856
rect 2706 711 3182 856
rect 3350 711 3826 856
rect 3994 711 4470 856
rect 4638 711 5114 856
rect 5282 711 6402 856
rect 6570 711 7046 856
rect 7214 711 7690 856
rect 7858 711 8334 856
rect 8502 711 8978 856
rect 9146 711 9622 856
rect 9790 711 10266 856
rect 10434 711 10910 856
rect 11078 711 12198 856
rect 12366 711 12842 856
rect 13010 711 13486 856
rect 13654 711 14130 856
rect 14298 711 14774 856
rect 14942 711 15418 856
rect 15586 711 16062 856
rect 16230 711 16706 856
rect 16874 711 17350 856
rect 17518 711 18638 856
rect 18806 711 19282 856
rect 19450 711 19926 856
rect 20094 711 20570 856
rect 20738 711 21214 856
rect 21382 711 21858 856
rect 22026 711 22502 856
rect 22670 711 23146 856
rect 23314 711 24434 856
rect 24602 711 25078 856
rect 25246 711 25722 856
rect 25890 711 26366 856
rect 26534 711 27010 856
rect 27178 711 27654 856
rect 27822 711 28298 856
rect 28466 711 28942 856
rect 29110 711 29586 856
rect 29754 711 30874 856
rect 31042 711 31518 856
rect 31686 711 32162 856
rect 32330 711 32806 856
rect 32974 711 33450 856
rect 33618 711 34094 856
rect 34262 711 34738 856
rect 34906 711 35382 856
rect 35550 711 36670 856
rect 36838 711 37314 856
rect 37482 711 37958 856
rect 38126 711 38602 856
rect 38770 711 39246 856
rect 39414 711 39890 856
rect 40058 711 40534 856
rect 40702 711 41178 856
rect 41346 711 41822 856
rect 41990 711 43110 856
rect 43278 711 43754 856
rect 43922 711 44398 856
rect 44566 711 45042 856
rect 45210 711 45686 856
rect 45854 711 46330 856
rect 46498 711 46974 856
rect 47142 711 47618 856
rect 47786 711 48906 856
rect 49074 711 49550 856
rect 49718 711 50194 856
rect 50362 711 50838 856
rect 51006 711 51482 856
rect 51650 711 52126 856
rect 52294 711 52770 856
rect 52938 711 53414 856
rect 53582 711 54058 856
rect 54226 711 55346 856
rect 55514 711 55990 856
rect 56158 711 56634 856
rect 56802 711 57278 856
rect 57446 711 57922 856
rect 58090 711 58566 856
rect 58734 711 59210 856
rect 59378 711 59854 856
rect 60022 711 61142 856
rect 61310 711 61786 856
rect 61954 711 62430 856
rect 62598 711 63074 856
rect 63242 711 63718 856
rect 63886 711 64362 856
rect 64530 711 65006 856
rect 65174 711 65650 856
rect 65818 711 66294 856
rect 66462 711 67582 856
rect 67750 711 68226 856
rect 68394 711 68870 856
rect 69038 711 69514 856
rect 69682 711 70158 856
rect 70326 711 70802 856
rect 70970 711 71446 856
rect 71614 711 72090 856
rect 72258 711 73378 856
rect 73546 711 74022 856
rect 74190 711 74666 856
rect 74834 711 75310 856
rect 75478 711 75954 856
rect 76122 711 76598 856
rect 76766 711 77242 856
rect 77410 711 77886 856
rect 78054 711 79174 856
rect 79342 711 79818 856
rect 79986 711 80462 856
rect 80630 711 81106 856
rect 81274 711 81750 856
rect 81918 711 82394 856
rect 82562 711 83038 856
rect 83206 711 83682 856
rect 83850 711 84326 856
rect 84494 711 85614 856
rect 85782 711 86258 856
rect 86426 711 86902 856
rect 87070 711 87546 856
rect 87714 711 88190 856
rect 88358 711 88834 856
rect 89002 711 89478 856
rect 89646 711 90122 856
rect 90290 711 91410 856
rect 91578 711 92054 856
rect 92222 711 92698 856
rect 92866 711 93342 856
rect 93510 711 93986 856
rect 94154 711 94630 856
rect 94798 711 95274 856
rect 95442 711 95918 856
rect 96086 711 96562 856
rect 96730 711 97850 856
rect 98018 711 98494 856
rect 98662 711 99138 856
rect 99306 711 99782 856
rect 99950 711 100426 856
rect 100594 711 101070 856
rect 101238 711 101714 856
rect 101882 711 102358 856
rect 102526 711 103646 856
rect 103814 711 104290 856
rect 104458 711 104934 856
rect 105102 711 105578 856
rect 105746 711 106222 856
rect 106390 711 106866 856
rect 107034 711 107510 856
rect 107678 711 108154 856
rect 108322 711 108798 856
rect 108966 711 110086 856
rect 110254 711 110730 856
rect 110898 711 111374 856
rect 111542 711 112018 856
rect 112186 711 112662 856
rect 112830 711 113306 856
rect 113474 711 113950 856
rect 114118 711 114594 856
rect 114762 711 115882 856
rect 116050 711 116526 856
rect 116694 711 117170 856
rect 117338 711 117814 856
rect 117982 711 118458 856
rect 118626 711 119102 856
rect 119270 711 119746 856
rect 119914 711 120390 856
rect 120558 711 121034 856
rect 121202 711 122322 856
rect 122490 711 122966 856
rect 123134 711 123610 856
rect 123778 711 124254 856
rect 124422 711 124898 856
rect 125066 711 125542 856
rect 125710 711 126186 856
rect 126354 711 126830 856
rect 126998 711 128118 856
rect 128286 711 128762 856
rect 128930 711 129406 856
rect 129574 711 130050 856
rect 130218 711 130694 856
rect 130862 711 131338 856
rect 131506 711 131982 856
rect 132150 711 132626 856
rect 132794 711 133270 856
rect 133438 711 134558 856
rect 134726 711 135202 856
rect 135370 711 135846 856
rect 136014 711 136490 856
rect 136658 711 137134 856
rect 137302 711 137778 856
rect 137946 711 138422 856
rect 138590 711 139066 856
rect 139234 711 140354 856
rect 140522 711 140998 856
rect 141166 711 141642 856
rect 141810 711 142286 856
rect 142454 711 142930 856
rect 143098 711 143574 856
rect 143742 711 144218 856
rect 144386 711 144862 856
rect 145030 711 145506 856
rect 145674 711 146794 856
rect 146962 711 147438 856
rect 147606 711 148082 856
rect 148250 711 148726 856
rect 148894 711 149370 856
rect 149538 711 150014 856
rect 150182 711 150658 856
rect 150826 711 151302 856
rect 151470 711 152590 856
rect 152758 711 153234 856
rect 153402 711 153878 856
rect 154046 711 154522 856
rect 154690 711 155166 856
rect 155334 711 155810 856
rect 155978 711 156454 856
rect 156622 711 157098 856
rect 157266 711 158386 856
rect 158554 711 159030 856
rect 159198 711 159674 856
rect 159842 711 160318 856
rect 160486 711 160962 856
rect 161130 711 161606 856
rect 161774 711 162250 856
rect 162418 711 162894 856
rect 163062 711 163538 856
rect 163706 711 164826 856
rect 164994 711 165470 856
rect 165638 711 166114 856
rect 166282 711 166758 856
rect 166926 711 167402 856
rect 167570 711 168046 856
rect 168214 711 168690 856
rect 168858 711 169334 856
rect 169502 711 170622 856
rect 170790 711 171266 856
rect 171434 711 171910 856
rect 172078 711 172554 856
rect 172722 711 173198 856
rect 173366 711 173842 856
rect 174010 711 174486 856
rect 174654 711 175130 856
rect 175298 711 175774 856
rect 175942 711 177062 856
rect 177230 711 177706 856
rect 177874 711 178350 856
rect 178518 711 178994 856
rect 179162 711 179638 856
rect 179806 711 180282 856
rect 180450 711 180926 856
rect 181094 711 181570 856
rect 181738 711 182858 856
rect 183026 711 183502 856
rect 183670 711 184146 856
rect 184314 711 184790 856
rect 184958 711 185434 856
rect 185602 711 186078 856
rect 186246 711 186722 856
rect 186890 711 187366 856
rect 187534 711 188010 856
rect 188178 711 189298 856
rect 189466 711 189942 856
rect 190110 711 190586 856
rect 190754 711 191230 856
rect 191398 711 191874 856
rect 192042 711 192518 856
rect 192686 711 193162 856
rect 193330 711 193806 856
rect 193974 711 195094 856
rect 195262 711 195738 856
rect 195906 711 196382 856
rect 196550 711 197026 856
rect 197194 711 197670 856
rect 197838 711 198314 856
rect 198482 711 198958 856
rect 199126 711 199602 856
rect 199770 711 200246 856
rect 200414 711 201534 856
rect 201702 711 202178 856
rect 202346 711 202822 856
rect 202990 711 203466 856
rect 203634 711 204110 856
rect 204278 711 204754 856
rect 204922 711 205398 856
rect 205566 711 206042 856
rect 206210 711 207330 856
rect 207498 711 207974 856
rect 208142 711 208618 856
rect 208786 711 209262 856
rect 209430 711 209906 856
rect 210074 711 210550 856
rect 210718 711 211194 856
rect 211362 711 211838 856
rect 212006 711 212482 856
rect 212650 711 213770 856
rect 213938 711 214414 856
rect 214582 711 215058 856
rect 215226 711 215702 856
rect 215870 711 216346 856
rect 216514 711 216990 856
rect 217158 711 217634 856
rect 217802 711 218278 856
rect 218446 711 219566 856
rect 219734 711 220210 856
rect 220378 711 220854 856
rect 221022 711 221498 856
rect 221666 711 222142 856
rect 222310 711 222786 856
rect 222954 711 223430 856
rect 223598 711 224074 856
rect 224242 711 224718 856
rect 224886 711 226006 856
rect 226174 711 226650 856
rect 226818 711 227294 856
rect 227462 711 227938 856
rect 228106 711 228582 856
rect 228750 711 229226 856
rect 229394 711 229870 856
rect 230038 711 230514 856
rect 230682 711 231802 856
rect 231970 711 232446 856
rect 232614 711 233090 856
rect 233258 711 233734 856
rect 233902 711 234378 856
rect 234546 711 235022 856
rect 235190 711 235666 856
rect 235834 711 236310 856
rect 236478 711 237598 856
rect 237766 711 238242 856
rect 238410 711 238886 856
rect 239054 711 239530 856
rect 239698 711 240174 856
rect 240342 711 240818 856
rect 240986 711 241462 856
rect 241630 711 242106 856
rect 242274 711 242750 856
rect 242918 711 244038 856
rect 244206 711 244682 856
rect 244850 711 245326 856
rect 245494 711 245970 856
rect 246138 711 246614 856
rect 246782 711 247258 856
rect 247426 711 247902 856
rect 248070 711 248546 856
rect 248714 711 249834 856
rect 250002 711 250478 856
rect 250646 711 251122 856
rect 251290 711 251766 856
rect 251934 711 252410 856
rect 252578 711 253054 856
rect 253222 711 253698 856
rect 253866 711 254342 856
rect 254510 711 254986 856
rect 255154 711 256274 856
rect 256442 711 256918 856
rect 257086 711 257562 856
rect 257730 711 258206 856
rect 258374 711 258850 856
rect 259018 711 259494 856
rect 259662 711 260138 856
rect 260306 711 260782 856
rect 260950 711 262070 856
rect 262238 711 262714 856
rect 262882 711 263358 856
rect 263526 711 264002 856
rect 264170 711 264646 856
rect 264814 711 265290 856
rect 265458 711 265934 856
rect 266102 711 266578 856
rect 266746 711 267222 856
rect 267390 711 268510 856
rect 268678 711 269154 856
rect 269322 711 269798 856
rect 269966 711 270442 856
rect 270610 711 271086 856
rect 271254 711 271730 856
rect 271898 711 272374 856
rect 272542 711 273018 856
rect 273186 711 274306 856
rect 274474 711 274950 856
rect 275118 711 275594 856
rect 275762 711 276238 856
rect 276406 711 276882 856
rect 277050 711 277526 856
rect 277694 711 278170 856
rect 278338 711 278814 856
rect 278982 711 279458 856
rect 279626 711 279660 856
<< metal3 >>
rect 279200 359728 280000 359848
rect 0 359048 800 359168
rect 279200 359048 280000 359168
rect 0 358368 800 358488
rect 279200 358368 280000 358488
rect 0 357688 800 357808
rect 279200 357688 280000 357808
rect 0 357008 800 357128
rect 279200 357008 280000 357128
rect 0 356328 800 356448
rect 279200 356328 280000 356448
rect 0 355648 800 355768
rect 279200 355648 280000 355768
rect 0 354968 800 355088
rect 279200 354968 280000 355088
rect 0 354288 800 354408
rect 279200 354288 280000 354408
rect 0 352928 800 353048
rect 279200 352928 280000 353048
rect 0 352248 800 352368
rect 279200 352248 280000 352368
rect 0 351568 800 351688
rect 279200 351568 280000 351688
rect 0 350888 800 351008
rect 279200 350888 280000 351008
rect 0 350208 800 350328
rect 279200 350208 280000 350328
rect 0 349528 800 349648
rect 279200 349528 280000 349648
rect 0 348848 800 348968
rect 279200 348848 280000 348968
rect 0 348168 800 348288
rect 279200 348168 280000 348288
rect 0 347488 800 347608
rect 279200 346808 280000 346928
rect 0 346128 800 346248
rect 279200 346128 280000 346248
rect 0 345448 800 345568
rect 279200 345448 280000 345568
rect 0 344768 800 344888
rect 279200 344768 280000 344888
rect 0 344088 800 344208
rect 279200 344088 280000 344208
rect 0 343408 800 343528
rect 279200 343408 280000 343528
rect 0 342728 800 342848
rect 279200 342728 280000 342848
rect 0 342048 800 342168
rect 279200 342048 280000 342168
rect 0 341368 800 341488
rect 279200 341368 280000 341488
rect 0 340008 800 340128
rect 279200 340008 280000 340128
rect 0 339328 800 339448
rect 279200 339328 280000 339448
rect 0 338648 800 338768
rect 279200 338648 280000 338768
rect 0 337968 800 338088
rect 279200 337968 280000 338088
rect 0 337288 800 337408
rect 279200 337288 280000 337408
rect 0 336608 800 336728
rect 279200 336608 280000 336728
rect 0 335928 800 336048
rect 279200 335928 280000 336048
rect 0 335248 800 335368
rect 279200 335248 280000 335368
rect 0 334568 800 334688
rect 279200 333888 280000 334008
rect 0 333208 800 333328
rect 279200 333208 280000 333328
rect 0 332528 800 332648
rect 279200 332528 280000 332648
rect 0 331848 800 331968
rect 279200 331848 280000 331968
rect 0 331168 800 331288
rect 279200 331168 280000 331288
rect 0 330488 800 330608
rect 279200 330488 280000 330608
rect 0 329808 800 329928
rect 279200 329808 280000 329928
rect 0 329128 800 329248
rect 279200 329128 280000 329248
rect 0 328448 800 328568
rect 279200 328448 280000 328568
rect 0 327088 800 327208
rect 279200 327088 280000 327208
rect 0 326408 800 326528
rect 279200 326408 280000 326528
rect 0 325728 800 325848
rect 279200 325728 280000 325848
rect 0 325048 800 325168
rect 279200 325048 280000 325168
rect 0 324368 800 324488
rect 279200 324368 280000 324488
rect 0 323688 800 323808
rect 279200 323688 280000 323808
rect 0 323008 800 323128
rect 279200 323008 280000 323128
rect 0 322328 800 322448
rect 279200 322328 280000 322448
rect 0 320968 800 321088
rect 279200 320968 280000 321088
rect 0 320288 800 320408
rect 279200 320288 280000 320408
rect 0 319608 800 319728
rect 279200 319608 280000 319728
rect 0 318928 800 319048
rect 279200 318928 280000 319048
rect 0 318248 800 318368
rect 279200 318248 280000 318368
rect 0 317568 800 317688
rect 279200 317568 280000 317688
rect 0 316888 800 317008
rect 279200 316888 280000 317008
rect 0 316208 800 316328
rect 279200 316208 280000 316328
rect 0 315528 800 315648
rect 279200 315528 280000 315648
rect 0 314168 800 314288
rect 279200 314168 280000 314288
rect 0 313488 800 313608
rect 279200 313488 280000 313608
rect 0 312808 800 312928
rect 279200 312808 280000 312928
rect 0 312128 800 312248
rect 279200 312128 280000 312248
rect 0 311448 800 311568
rect 279200 311448 280000 311568
rect 0 310768 800 310888
rect 279200 310768 280000 310888
rect 0 310088 800 310208
rect 279200 310088 280000 310208
rect 0 309408 800 309528
rect 279200 309408 280000 309528
rect 0 308048 800 308168
rect 279200 308048 280000 308168
rect 0 307368 800 307488
rect 279200 307368 280000 307488
rect 0 306688 800 306808
rect 279200 306688 280000 306808
rect 0 306008 800 306128
rect 279200 306008 280000 306128
rect 0 305328 800 305448
rect 279200 305328 280000 305448
rect 0 304648 800 304768
rect 279200 304648 280000 304768
rect 0 303968 800 304088
rect 279200 303968 280000 304088
rect 0 303288 800 303408
rect 279200 303288 280000 303408
rect 0 302608 800 302728
rect 279200 302608 280000 302728
rect 0 301248 800 301368
rect 279200 301248 280000 301368
rect 0 300568 800 300688
rect 279200 300568 280000 300688
rect 0 299888 800 300008
rect 279200 299888 280000 300008
rect 0 299208 800 299328
rect 279200 299208 280000 299328
rect 0 298528 800 298648
rect 279200 298528 280000 298648
rect 0 297848 800 297968
rect 279200 297848 280000 297968
rect 0 297168 800 297288
rect 279200 297168 280000 297288
rect 0 296488 800 296608
rect 279200 296488 280000 296608
rect 0 295128 800 295248
rect 279200 295128 280000 295248
rect 0 294448 800 294568
rect 279200 294448 280000 294568
rect 0 293768 800 293888
rect 279200 293768 280000 293888
rect 0 293088 800 293208
rect 279200 293088 280000 293208
rect 0 292408 800 292528
rect 279200 292408 280000 292528
rect 0 291728 800 291848
rect 279200 291728 280000 291848
rect 0 291048 800 291168
rect 279200 291048 280000 291168
rect 0 290368 800 290488
rect 279200 290368 280000 290488
rect 0 289688 800 289808
rect 279200 289688 280000 289808
rect 0 288328 800 288448
rect 279200 288328 280000 288448
rect 0 287648 800 287768
rect 279200 287648 280000 287768
rect 0 286968 800 287088
rect 279200 286968 280000 287088
rect 0 286288 800 286408
rect 279200 286288 280000 286408
rect 0 285608 800 285728
rect 279200 285608 280000 285728
rect 0 284928 800 285048
rect 279200 284928 280000 285048
rect 0 284248 800 284368
rect 279200 284248 280000 284368
rect 0 283568 800 283688
rect 279200 283568 280000 283688
rect 0 282208 800 282328
rect 279200 282208 280000 282328
rect 0 281528 800 281648
rect 279200 281528 280000 281648
rect 0 280848 800 280968
rect 279200 280848 280000 280968
rect 0 280168 800 280288
rect 279200 280168 280000 280288
rect 0 279488 800 279608
rect 279200 279488 280000 279608
rect 0 278808 800 278928
rect 279200 278808 280000 278928
rect 0 278128 800 278248
rect 279200 278128 280000 278248
rect 0 277448 800 277568
rect 279200 277448 280000 277568
rect 0 276768 800 276888
rect 279200 276088 280000 276208
rect 0 275408 800 275528
rect 279200 275408 280000 275528
rect 0 274728 800 274848
rect 279200 274728 280000 274848
rect 0 274048 800 274168
rect 279200 274048 280000 274168
rect 0 273368 800 273488
rect 279200 273368 280000 273488
rect 0 272688 800 272808
rect 279200 272688 280000 272808
rect 0 272008 800 272128
rect 279200 272008 280000 272128
rect 0 271328 800 271448
rect 279200 271328 280000 271448
rect 0 270648 800 270768
rect 279200 270648 280000 270768
rect 0 269288 800 269408
rect 279200 269288 280000 269408
rect 0 268608 800 268728
rect 279200 268608 280000 268728
rect 0 267928 800 268048
rect 279200 267928 280000 268048
rect 0 267248 800 267368
rect 279200 267248 280000 267368
rect 0 266568 800 266688
rect 279200 266568 280000 266688
rect 0 265888 800 266008
rect 279200 265888 280000 266008
rect 0 265208 800 265328
rect 279200 265208 280000 265328
rect 0 264528 800 264648
rect 279200 264528 280000 264648
rect 0 263848 800 263968
rect 279200 263168 280000 263288
rect 0 262488 800 262608
rect 279200 262488 280000 262608
rect 0 261808 800 261928
rect 279200 261808 280000 261928
rect 0 261128 800 261248
rect 279200 261128 280000 261248
rect 0 260448 800 260568
rect 279200 260448 280000 260568
rect 0 259768 800 259888
rect 279200 259768 280000 259888
rect 0 259088 800 259208
rect 279200 259088 280000 259208
rect 0 258408 800 258528
rect 279200 258408 280000 258528
rect 0 257728 800 257848
rect 279200 257728 280000 257848
rect 0 256368 800 256488
rect 279200 256368 280000 256488
rect 0 255688 800 255808
rect 279200 255688 280000 255808
rect 0 255008 800 255128
rect 279200 255008 280000 255128
rect 0 254328 800 254448
rect 279200 254328 280000 254448
rect 0 253648 800 253768
rect 279200 253648 280000 253768
rect 0 252968 800 253088
rect 279200 252968 280000 253088
rect 0 252288 800 252408
rect 279200 252288 280000 252408
rect 0 251608 800 251728
rect 279200 251608 280000 251728
rect 0 250928 800 251048
rect 279200 250248 280000 250368
rect 0 249568 800 249688
rect 279200 249568 280000 249688
rect 0 248888 800 249008
rect 279200 248888 280000 249008
rect 0 248208 800 248328
rect 279200 248208 280000 248328
rect 0 247528 800 247648
rect 279200 247528 280000 247648
rect 0 246848 800 246968
rect 279200 246848 280000 246968
rect 0 246168 800 246288
rect 279200 246168 280000 246288
rect 0 245488 800 245608
rect 279200 245488 280000 245608
rect 0 244808 800 244928
rect 279200 244808 280000 244928
rect 0 243448 800 243568
rect 279200 243448 280000 243568
rect 0 242768 800 242888
rect 279200 242768 280000 242888
rect 0 242088 800 242208
rect 279200 242088 280000 242208
rect 0 241408 800 241528
rect 279200 241408 280000 241528
rect 0 240728 800 240848
rect 279200 240728 280000 240848
rect 0 240048 800 240168
rect 279200 240048 280000 240168
rect 0 239368 800 239488
rect 279200 239368 280000 239488
rect 0 238688 800 238808
rect 279200 238688 280000 238808
rect 0 237328 800 237448
rect 279200 237328 280000 237448
rect 0 236648 800 236768
rect 279200 236648 280000 236768
rect 0 235968 800 236088
rect 279200 235968 280000 236088
rect 0 235288 800 235408
rect 279200 235288 280000 235408
rect 0 234608 800 234728
rect 279200 234608 280000 234728
rect 0 233928 800 234048
rect 279200 233928 280000 234048
rect 0 233248 800 233368
rect 279200 233248 280000 233368
rect 0 232568 800 232688
rect 279200 232568 280000 232688
rect 0 231888 800 232008
rect 279200 231888 280000 232008
rect 0 230528 800 230648
rect 279200 230528 280000 230648
rect 0 229848 800 229968
rect 279200 229848 280000 229968
rect 0 229168 800 229288
rect 279200 229168 280000 229288
rect 0 228488 800 228608
rect 279200 228488 280000 228608
rect 0 227808 800 227928
rect 279200 227808 280000 227928
rect 0 227128 800 227248
rect 279200 227128 280000 227248
rect 0 226448 800 226568
rect 279200 226448 280000 226568
rect 0 225768 800 225888
rect 279200 225768 280000 225888
rect 0 224408 800 224528
rect 279200 224408 280000 224528
rect 0 223728 800 223848
rect 279200 223728 280000 223848
rect 0 223048 800 223168
rect 279200 223048 280000 223168
rect 0 222368 800 222488
rect 279200 222368 280000 222488
rect 0 221688 800 221808
rect 279200 221688 280000 221808
rect 0 221008 800 221128
rect 279200 221008 280000 221128
rect 0 220328 800 220448
rect 279200 220328 280000 220448
rect 0 219648 800 219768
rect 279200 219648 280000 219768
rect 0 218968 800 219088
rect 279200 218968 280000 219088
rect 0 217608 800 217728
rect 279200 217608 280000 217728
rect 0 216928 800 217048
rect 279200 216928 280000 217048
rect 0 216248 800 216368
rect 279200 216248 280000 216368
rect 0 215568 800 215688
rect 279200 215568 280000 215688
rect 0 214888 800 215008
rect 279200 214888 280000 215008
rect 0 214208 800 214328
rect 279200 214208 280000 214328
rect 0 213528 800 213648
rect 279200 213528 280000 213648
rect 0 212848 800 212968
rect 279200 212848 280000 212968
rect 0 211488 800 211608
rect 279200 211488 280000 211608
rect 0 210808 800 210928
rect 279200 210808 280000 210928
rect 0 210128 800 210248
rect 279200 210128 280000 210248
rect 0 209448 800 209568
rect 279200 209448 280000 209568
rect 0 208768 800 208888
rect 279200 208768 280000 208888
rect 0 208088 800 208208
rect 279200 208088 280000 208208
rect 0 207408 800 207528
rect 279200 207408 280000 207528
rect 0 206728 800 206848
rect 279200 206728 280000 206848
rect 0 206048 800 206168
rect 279200 206048 280000 206168
rect 0 204688 800 204808
rect 279200 204688 280000 204808
rect 0 204008 800 204128
rect 279200 204008 280000 204128
rect 0 203328 800 203448
rect 279200 203328 280000 203448
rect 0 202648 800 202768
rect 279200 202648 280000 202768
rect 0 201968 800 202088
rect 279200 201968 280000 202088
rect 0 201288 800 201408
rect 279200 201288 280000 201408
rect 0 200608 800 200728
rect 279200 200608 280000 200728
rect 0 199928 800 200048
rect 279200 199928 280000 200048
rect 0 198568 800 198688
rect 279200 198568 280000 198688
rect 0 197888 800 198008
rect 279200 197888 280000 198008
rect 0 197208 800 197328
rect 279200 197208 280000 197328
rect 0 196528 800 196648
rect 279200 196528 280000 196648
rect 0 195848 800 195968
rect 279200 195848 280000 195968
rect 0 195168 800 195288
rect 279200 195168 280000 195288
rect 0 194488 800 194608
rect 279200 194488 280000 194608
rect 0 193808 800 193928
rect 279200 193808 280000 193928
rect 0 193128 800 193248
rect 279200 192448 280000 192568
rect 0 191768 800 191888
rect 279200 191768 280000 191888
rect 0 191088 800 191208
rect 279200 191088 280000 191208
rect 0 190408 800 190528
rect 279200 190408 280000 190528
rect 0 189728 800 189848
rect 279200 189728 280000 189848
rect 0 189048 800 189168
rect 279200 189048 280000 189168
rect 0 188368 800 188488
rect 279200 188368 280000 188488
rect 0 187688 800 187808
rect 279200 187688 280000 187808
rect 0 187008 800 187128
rect 279200 187008 280000 187128
rect 0 185648 800 185768
rect 279200 185648 280000 185768
rect 0 184968 800 185088
rect 279200 184968 280000 185088
rect 0 184288 800 184408
rect 279200 184288 280000 184408
rect 0 183608 800 183728
rect 279200 183608 280000 183728
rect 0 182928 800 183048
rect 279200 182928 280000 183048
rect 0 182248 800 182368
rect 279200 182248 280000 182368
rect 0 181568 800 181688
rect 279200 181568 280000 181688
rect 0 180888 800 181008
rect 279200 180888 280000 181008
rect 0 180208 800 180328
rect 279200 179528 280000 179648
rect 0 178848 800 178968
rect 279200 178848 280000 178968
rect 0 178168 800 178288
rect 279200 178168 280000 178288
rect 0 177488 800 177608
rect 279200 177488 280000 177608
rect 0 176808 800 176928
rect 279200 176808 280000 176928
rect 0 176128 800 176248
rect 279200 176128 280000 176248
rect 0 175448 800 175568
rect 279200 175448 280000 175568
rect 0 174768 800 174888
rect 279200 174768 280000 174888
rect 0 174088 800 174208
rect 279200 174088 280000 174208
rect 0 172728 800 172848
rect 279200 172728 280000 172848
rect 0 172048 800 172168
rect 279200 172048 280000 172168
rect 0 171368 800 171488
rect 279200 171368 280000 171488
rect 0 170688 800 170808
rect 279200 170688 280000 170808
rect 0 170008 800 170128
rect 279200 170008 280000 170128
rect 0 169328 800 169448
rect 279200 169328 280000 169448
rect 0 168648 800 168768
rect 279200 168648 280000 168768
rect 0 167968 800 168088
rect 279200 167968 280000 168088
rect 0 167288 800 167408
rect 279200 166608 280000 166728
rect 0 165928 800 166048
rect 279200 165928 280000 166048
rect 0 165248 800 165368
rect 279200 165248 280000 165368
rect 0 164568 800 164688
rect 279200 164568 280000 164688
rect 0 163888 800 164008
rect 279200 163888 280000 164008
rect 0 163208 800 163328
rect 279200 163208 280000 163328
rect 0 162528 800 162648
rect 279200 162528 280000 162648
rect 0 161848 800 161968
rect 279200 161848 280000 161968
rect 0 161168 800 161288
rect 279200 161168 280000 161288
rect 0 159808 800 159928
rect 279200 159808 280000 159928
rect 0 159128 800 159248
rect 279200 159128 280000 159248
rect 0 158448 800 158568
rect 279200 158448 280000 158568
rect 0 157768 800 157888
rect 279200 157768 280000 157888
rect 0 157088 800 157208
rect 279200 157088 280000 157208
rect 0 156408 800 156528
rect 279200 156408 280000 156528
rect 0 155728 800 155848
rect 279200 155728 280000 155848
rect 0 155048 800 155168
rect 279200 155048 280000 155168
rect 0 153688 800 153808
rect 279200 153688 280000 153808
rect 0 153008 800 153128
rect 279200 153008 280000 153128
rect 0 152328 800 152448
rect 279200 152328 280000 152448
rect 0 151648 800 151768
rect 279200 151648 280000 151768
rect 0 150968 800 151088
rect 279200 150968 280000 151088
rect 0 150288 800 150408
rect 279200 150288 280000 150408
rect 0 149608 800 149728
rect 279200 149608 280000 149728
rect 0 148928 800 149048
rect 279200 148928 280000 149048
rect 0 148248 800 148368
rect 279200 148248 280000 148368
rect 0 146888 800 147008
rect 279200 146888 280000 147008
rect 0 146208 800 146328
rect 279200 146208 280000 146328
rect 0 145528 800 145648
rect 279200 145528 280000 145648
rect 0 144848 800 144968
rect 279200 144848 280000 144968
rect 0 144168 800 144288
rect 279200 144168 280000 144288
rect 0 143488 800 143608
rect 279200 143488 280000 143608
rect 0 142808 800 142928
rect 279200 142808 280000 142928
rect 0 142128 800 142248
rect 279200 142128 280000 142248
rect 0 140768 800 140888
rect 279200 140768 280000 140888
rect 0 140088 800 140208
rect 279200 140088 280000 140208
rect 0 139408 800 139528
rect 279200 139408 280000 139528
rect 0 138728 800 138848
rect 279200 138728 280000 138848
rect 0 138048 800 138168
rect 279200 138048 280000 138168
rect 0 137368 800 137488
rect 279200 137368 280000 137488
rect 0 136688 800 136808
rect 279200 136688 280000 136808
rect 0 136008 800 136128
rect 279200 136008 280000 136128
rect 0 135328 800 135448
rect 279200 135328 280000 135448
rect 0 133968 800 134088
rect 279200 133968 280000 134088
rect 0 133288 800 133408
rect 279200 133288 280000 133408
rect 0 132608 800 132728
rect 279200 132608 280000 132728
rect 0 131928 800 132048
rect 279200 131928 280000 132048
rect 0 131248 800 131368
rect 279200 131248 280000 131368
rect 0 130568 800 130688
rect 279200 130568 280000 130688
rect 0 129888 800 130008
rect 279200 129888 280000 130008
rect 0 129208 800 129328
rect 279200 129208 280000 129328
rect 0 127848 800 127968
rect 279200 127848 280000 127968
rect 0 127168 800 127288
rect 279200 127168 280000 127288
rect 0 126488 800 126608
rect 279200 126488 280000 126608
rect 0 125808 800 125928
rect 279200 125808 280000 125928
rect 0 125128 800 125248
rect 279200 125128 280000 125248
rect 0 124448 800 124568
rect 279200 124448 280000 124568
rect 0 123768 800 123888
rect 279200 123768 280000 123888
rect 0 123088 800 123208
rect 279200 123088 280000 123208
rect 0 122408 800 122528
rect 279200 122408 280000 122528
rect 0 121048 800 121168
rect 279200 121048 280000 121168
rect 0 120368 800 120488
rect 279200 120368 280000 120488
rect 0 119688 800 119808
rect 279200 119688 280000 119808
rect 0 119008 800 119128
rect 279200 119008 280000 119128
rect 0 118328 800 118448
rect 279200 118328 280000 118448
rect 0 117648 800 117768
rect 279200 117648 280000 117768
rect 0 116968 800 117088
rect 279200 116968 280000 117088
rect 0 116288 800 116408
rect 279200 116288 280000 116408
rect 0 114928 800 115048
rect 279200 114928 280000 115048
rect 0 114248 800 114368
rect 279200 114248 280000 114368
rect 0 113568 800 113688
rect 279200 113568 280000 113688
rect 0 112888 800 113008
rect 279200 112888 280000 113008
rect 0 112208 800 112328
rect 279200 112208 280000 112328
rect 0 111528 800 111648
rect 279200 111528 280000 111648
rect 0 110848 800 110968
rect 279200 110848 280000 110968
rect 0 110168 800 110288
rect 279200 110168 280000 110288
rect 0 109488 800 109608
rect 279200 108808 280000 108928
rect 0 108128 800 108248
rect 279200 108128 280000 108248
rect 0 107448 800 107568
rect 279200 107448 280000 107568
rect 0 106768 800 106888
rect 279200 106768 280000 106888
rect 0 106088 800 106208
rect 279200 106088 280000 106208
rect 0 105408 800 105528
rect 279200 105408 280000 105528
rect 0 104728 800 104848
rect 279200 104728 280000 104848
rect 0 104048 800 104168
rect 279200 104048 280000 104168
rect 0 103368 800 103488
rect 279200 103368 280000 103488
rect 0 102008 800 102128
rect 279200 102008 280000 102128
rect 0 101328 800 101448
rect 279200 101328 280000 101448
rect 0 100648 800 100768
rect 279200 100648 280000 100768
rect 0 99968 800 100088
rect 279200 99968 280000 100088
rect 0 99288 800 99408
rect 279200 99288 280000 99408
rect 0 98608 800 98728
rect 279200 98608 280000 98728
rect 0 97928 800 98048
rect 279200 97928 280000 98048
rect 0 97248 800 97368
rect 279200 97248 280000 97368
rect 0 96568 800 96688
rect 279200 95888 280000 96008
rect 0 95208 800 95328
rect 279200 95208 280000 95328
rect 0 94528 800 94648
rect 279200 94528 280000 94648
rect 0 93848 800 93968
rect 279200 93848 280000 93968
rect 0 93168 800 93288
rect 279200 93168 280000 93288
rect 0 92488 800 92608
rect 279200 92488 280000 92608
rect 0 91808 800 91928
rect 279200 91808 280000 91928
rect 0 91128 800 91248
rect 279200 91128 280000 91248
rect 0 90448 800 90568
rect 279200 90448 280000 90568
rect 0 89088 800 89208
rect 279200 89088 280000 89208
rect 0 88408 800 88528
rect 279200 88408 280000 88528
rect 0 87728 800 87848
rect 279200 87728 280000 87848
rect 0 87048 800 87168
rect 279200 87048 280000 87168
rect 0 86368 800 86488
rect 279200 86368 280000 86488
rect 0 85688 800 85808
rect 279200 85688 280000 85808
rect 0 85008 800 85128
rect 279200 85008 280000 85128
rect 0 84328 800 84448
rect 279200 84328 280000 84448
rect 0 83648 800 83768
rect 279200 82968 280000 83088
rect 0 82288 800 82408
rect 279200 82288 280000 82408
rect 0 81608 800 81728
rect 279200 81608 280000 81728
rect 0 80928 800 81048
rect 279200 80928 280000 81048
rect 0 80248 800 80368
rect 279200 80248 280000 80368
rect 0 79568 800 79688
rect 279200 79568 280000 79688
rect 0 78888 800 79008
rect 279200 78888 280000 79008
rect 0 78208 800 78328
rect 279200 78208 280000 78328
rect 0 77528 800 77648
rect 279200 77528 280000 77648
rect 0 76168 800 76288
rect 279200 76168 280000 76288
rect 0 75488 800 75608
rect 279200 75488 280000 75608
rect 0 74808 800 74928
rect 279200 74808 280000 74928
rect 0 74128 800 74248
rect 279200 74128 280000 74248
rect 0 73448 800 73568
rect 279200 73448 280000 73568
rect 0 72768 800 72888
rect 279200 72768 280000 72888
rect 0 72088 800 72208
rect 279200 72088 280000 72208
rect 0 71408 800 71528
rect 279200 71408 280000 71528
rect 0 70048 800 70168
rect 279200 70048 280000 70168
rect 0 69368 800 69488
rect 279200 69368 280000 69488
rect 0 68688 800 68808
rect 279200 68688 280000 68808
rect 0 68008 800 68128
rect 279200 68008 280000 68128
rect 0 67328 800 67448
rect 279200 67328 280000 67448
rect 0 66648 800 66768
rect 279200 66648 280000 66768
rect 0 65968 800 66088
rect 279200 65968 280000 66088
rect 0 65288 800 65408
rect 279200 65288 280000 65408
rect 0 64608 800 64728
rect 279200 64608 280000 64728
rect 0 63248 800 63368
rect 279200 63248 280000 63368
rect 0 62568 800 62688
rect 279200 62568 280000 62688
rect 0 61888 800 62008
rect 279200 61888 280000 62008
rect 0 61208 800 61328
rect 279200 61208 280000 61328
rect 0 60528 800 60648
rect 279200 60528 280000 60648
rect 0 59848 800 59968
rect 279200 59848 280000 59968
rect 0 59168 800 59288
rect 279200 59168 280000 59288
rect 0 58488 800 58608
rect 279200 58488 280000 58608
rect 0 57128 800 57248
rect 279200 57128 280000 57248
rect 0 56448 800 56568
rect 279200 56448 280000 56568
rect 0 55768 800 55888
rect 279200 55768 280000 55888
rect 0 55088 800 55208
rect 279200 55088 280000 55208
rect 0 54408 800 54528
rect 279200 54408 280000 54528
rect 0 53728 800 53848
rect 279200 53728 280000 53848
rect 0 53048 800 53168
rect 279200 53048 280000 53168
rect 0 52368 800 52488
rect 279200 52368 280000 52488
rect 0 51688 800 51808
rect 279200 51688 280000 51808
rect 0 50328 800 50448
rect 279200 50328 280000 50448
rect 0 49648 800 49768
rect 279200 49648 280000 49768
rect 0 48968 800 49088
rect 279200 48968 280000 49088
rect 0 48288 800 48408
rect 279200 48288 280000 48408
rect 0 47608 800 47728
rect 279200 47608 280000 47728
rect 0 46928 800 47048
rect 279200 46928 280000 47048
rect 0 46248 800 46368
rect 279200 46248 280000 46368
rect 0 45568 800 45688
rect 279200 45568 280000 45688
rect 0 44208 800 44328
rect 279200 44208 280000 44328
rect 0 43528 800 43648
rect 279200 43528 280000 43648
rect 0 42848 800 42968
rect 279200 42848 280000 42968
rect 0 42168 800 42288
rect 279200 42168 280000 42288
rect 0 41488 800 41608
rect 279200 41488 280000 41608
rect 0 40808 800 40928
rect 279200 40808 280000 40928
rect 0 40128 800 40248
rect 279200 40128 280000 40248
rect 0 39448 800 39568
rect 279200 39448 280000 39568
rect 0 38768 800 38888
rect 279200 38768 280000 38888
rect 0 37408 800 37528
rect 279200 37408 280000 37528
rect 0 36728 800 36848
rect 279200 36728 280000 36848
rect 0 36048 800 36168
rect 279200 36048 280000 36168
rect 0 35368 800 35488
rect 279200 35368 280000 35488
rect 0 34688 800 34808
rect 279200 34688 280000 34808
rect 0 34008 800 34128
rect 279200 34008 280000 34128
rect 0 33328 800 33448
rect 279200 33328 280000 33448
rect 0 32648 800 32768
rect 279200 32648 280000 32768
rect 0 31288 800 31408
rect 279200 31288 280000 31408
rect 0 30608 800 30728
rect 279200 30608 280000 30728
rect 0 29928 800 30048
rect 279200 29928 280000 30048
rect 0 29248 800 29368
rect 279200 29248 280000 29368
rect 0 28568 800 28688
rect 279200 28568 280000 28688
rect 0 27888 800 28008
rect 279200 27888 280000 28008
rect 0 27208 800 27328
rect 279200 27208 280000 27328
rect 0 26528 800 26648
rect 279200 26528 280000 26648
rect 0 25848 800 25968
rect 279200 25168 280000 25288
rect 0 24488 800 24608
rect 279200 24488 280000 24608
rect 0 23808 800 23928
rect 279200 23808 280000 23928
rect 0 23128 800 23248
rect 279200 23128 280000 23248
rect 0 22448 800 22568
rect 279200 22448 280000 22568
rect 0 21768 800 21888
rect 279200 21768 280000 21888
rect 0 21088 800 21208
rect 279200 21088 280000 21208
rect 0 20408 800 20528
rect 279200 20408 280000 20528
rect 0 19728 800 19848
rect 279200 19728 280000 19848
rect 0 18368 800 18488
rect 279200 18368 280000 18488
rect 0 17688 800 17808
rect 279200 17688 280000 17808
rect 0 17008 800 17128
rect 279200 17008 280000 17128
rect 0 16328 800 16448
rect 279200 16328 280000 16448
rect 0 15648 800 15768
rect 279200 15648 280000 15768
rect 0 14968 800 15088
rect 279200 14968 280000 15088
rect 0 14288 800 14408
rect 279200 14288 280000 14408
rect 0 13608 800 13728
rect 279200 13608 280000 13728
rect 0 12928 800 13048
rect 279200 12248 280000 12368
rect 0 11568 800 11688
rect 279200 11568 280000 11688
rect 0 10888 800 11008
rect 279200 10888 280000 11008
rect 0 10208 800 10328
rect 279200 10208 280000 10328
rect 0 9528 800 9648
rect 279200 9528 280000 9648
rect 0 8848 800 8968
rect 279200 8848 280000 8968
rect 0 8168 800 8288
rect 279200 8168 280000 8288
rect 0 7488 800 7608
rect 279200 7488 280000 7608
rect 0 6808 800 6928
rect 279200 6808 280000 6928
rect 0 5448 800 5568
rect 279200 5448 280000 5568
rect 0 4768 800 4888
rect 279200 4768 280000 4888
rect 0 4088 800 4208
rect 279200 4088 280000 4208
rect 0 3408 800 3528
rect 279200 3408 280000 3528
rect 0 2728 800 2848
rect 279200 2728 280000 2848
rect 0 2048 800 2168
rect 279200 2048 280000 2168
rect 0 1368 800 1488
rect 279200 1368 280000 1488
rect 0 688 800 808
rect 279200 688 280000 808
<< obsm3 >>
rect 880 358968 279120 359141
rect 565 358568 279575 358968
rect 880 358288 279120 358568
rect 565 357888 279575 358288
rect 880 357608 279120 357888
rect 565 357208 279575 357608
rect 880 356928 279120 357208
rect 565 356528 279575 356928
rect 880 356248 279120 356528
rect 565 355848 279575 356248
rect 880 355568 279120 355848
rect 565 355168 279575 355568
rect 880 354888 279120 355168
rect 565 354488 279575 354888
rect 880 354208 279120 354488
rect 565 353128 279575 354208
rect 880 352848 279120 353128
rect 565 352448 279575 352848
rect 880 352168 279120 352448
rect 565 351768 279575 352168
rect 880 351488 279120 351768
rect 565 351088 279575 351488
rect 880 350808 279120 351088
rect 565 350408 279575 350808
rect 880 350128 279120 350408
rect 565 349728 279575 350128
rect 880 349448 279120 349728
rect 565 349048 279575 349448
rect 880 348768 279120 349048
rect 565 348368 279575 348768
rect 880 348088 279120 348368
rect 565 347688 279575 348088
rect 880 347408 279575 347688
rect 565 347008 279575 347408
rect 565 346728 279120 347008
rect 565 346328 279575 346728
rect 880 346048 279120 346328
rect 565 345648 279575 346048
rect 880 345368 279120 345648
rect 565 344968 279575 345368
rect 880 344688 279120 344968
rect 565 344288 279575 344688
rect 880 344008 279120 344288
rect 565 343608 279575 344008
rect 880 343328 279120 343608
rect 565 342928 279575 343328
rect 880 342648 279120 342928
rect 565 342248 279575 342648
rect 880 341968 279120 342248
rect 565 341568 279575 341968
rect 880 341288 279120 341568
rect 565 340208 279575 341288
rect 880 339928 279120 340208
rect 565 339528 279575 339928
rect 880 339248 279120 339528
rect 565 338848 279575 339248
rect 880 338568 279120 338848
rect 565 338168 279575 338568
rect 880 337888 279120 338168
rect 565 337488 279575 337888
rect 880 337208 279120 337488
rect 565 336808 279575 337208
rect 880 336528 279120 336808
rect 565 336128 279575 336528
rect 880 335848 279120 336128
rect 565 335448 279575 335848
rect 880 335168 279120 335448
rect 565 334768 279575 335168
rect 880 334488 279575 334768
rect 565 334088 279575 334488
rect 565 333808 279120 334088
rect 565 333408 279575 333808
rect 880 333128 279120 333408
rect 565 332728 279575 333128
rect 880 332448 279120 332728
rect 565 332048 279575 332448
rect 880 331768 279120 332048
rect 565 331368 279575 331768
rect 880 331088 279120 331368
rect 565 330688 279575 331088
rect 880 330408 279120 330688
rect 565 330008 279575 330408
rect 880 329728 279120 330008
rect 565 329328 279575 329728
rect 880 329048 279120 329328
rect 565 328648 279575 329048
rect 880 328368 279120 328648
rect 565 327288 279575 328368
rect 880 327008 279120 327288
rect 565 326608 279575 327008
rect 880 326328 279120 326608
rect 565 325928 279575 326328
rect 880 325648 279120 325928
rect 565 325248 279575 325648
rect 880 324968 279120 325248
rect 565 324568 279575 324968
rect 880 324288 279120 324568
rect 565 323888 279575 324288
rect 880 323608 279120 323888
rect 565 323208 279575 323608
rect 880 322928 279120 323208
rect 565 322528 279575 322928
rect 880 322248 279120 322528
rect 565 321168 279575 322248
rect 880 320888 279120 321168
rect 565 320488 279575 320888
rect 880 320208 279120 320488
rect 565 319808 279575 320208
rect 880 319528 279120 319808
rect 565 319128 279575 319528
rect 880 318848 279120 319128
rect 565 318448 279575 318848
rect 880 318168 279120 318448
rect 565 317768 279575 318168
rect 880 317488 279120 317768
rect 565 317088 279575 317488
rect 880 316808 279120 317088
rect 565 316408 279575 316808
rect 880 316128 279120 316408
rect 565 315728 279575 316128
rect 880 315448 279120 315728
rect 565 314368 279575 315448
rect 880 314088 279120 314368
rect 565 313688 279575 314088
rect 880 313408 279120 313688
rect 565 313008 279575 313408
rect 880 312728 279120 313008
rect 565 312328 279575 312728
rect 880 312048 279120 312328
rect 565 311648 279575 312048
rect 880 311368 279120 311648
rect 565 310968 279575 311368
rect 880 310688 279120 310968
rect 565 310288 279575 310688
rect 880 310008 279120 310288
rect 565 309608 279575 310008
rect 880 309328 279120 309608
rect 565 308248 279575 309328
rect 880 307968 279120 308248
rect 565 307568 279575 307968
rect 880 307288 279120 307568
rect 565 306888 279575 307288
rect 880 306608 279120 306888
rect 565 306208 279575 306608
rect 880 305928 279120 306208
rect 565 305528 279575 305928
rect 880 305248 279120 305528
rect 565 304848 279575 305248
rect 880 304568 279120 304848
rect 565 304168 279575 304568
rect 880 303888 279120 304168
rect 565 303488 279575 303888
rect 880 303208 279120 303488
rect 565 302808 279575 303208
rect 880 302528 279120 302808
rect 565 301448 279575 302528
rect 880 301168 279120 301448
rect 565 300768 279575 301168
rect 880 300488 279120 300768
rect 565 300088 279575 300488
rect 880 299808 279120 300088
rect 565 299408 279575 299808
rect 880 299128 279120 299408
rect 565 298728 279575 299128
rect 880 298448 279120 298728
rect 565 298048 279575 298448
rect 880 297768 279120 298048
rect 565 297368 279575 297768
rect 880 297088 279120 297368
rect 565 296688 279575 297088
rect 880 296408 279120 296688
rect 565 295328 279575 296408
rect 880 295048 279120 295328
rect 565 294648 279575 295048
rect 880 294368 279120 294648
rect 565 293968 279575 294368
rect 880 293688 279120 293968
rect 565 293288 279575 293688
rect 880 293008 279120 293288
rect 565 292608 279575 293008
rect 880 292328 279120 292608
rect 565 291928 279575 292328
rect 880 291648 279120 291928
rect 565 291248 279575 291648
rect 880 290968 279120 291248
rect 565 290568 279575 290968
rect 880 290288 279120 290568
rect 565 289888 279575 290288
rect 880 289608 279120 289888
rect 565 288528 279575 289608
rect 880 288248 279120 288528
rect 565 287848 279575 288248
rect 880 287568 279120 287848
rect 565 287168 279575 287568
rect 880 286888 279120 287168
rect 565 286488 279575 286888
rect 880 286208 279120 286488
rect 565 285808 279575 286208
rect 880 285528 279120 285808
rect 565 285128 279575 285528
rect 880 284848 279120 285128
rect 565 284448 279575 284848
rect 880 284168 279120 284448
rect 565 283768 279575 284168
rect 880 283488 279120 283768
rect 565 282408 279575 283488
rect 880 282128 279120 282408
rect 565 281728 279575 282128
rect 880 281448 279120 281728
rect 565 281048 279575 281448
rect 880 280768 279120 281048
rect 565 280368 279575 280768
rect 880 280088 279120 280368
rect 565 279688 279575 280088
rect 880 279408 279120 279688
rect 565 279008 279575 279408
rect 880 278728 279120 279008
rect 565 278328 279575 278728
rect 880 278048 279120 278328
rect 565 277648 279575 278048
rect 880 277368 279120 277648
rect 565 276968 279575 277368
rect 880 276688 279575 276968
rect 565 276288 279575 276688
rect 565 276008 279120 276288
rect 565 275608 279575 276008
rect 880 275328 279120 275608
rect 565 274928 279575 275328
rect 880 274648 279120 274928
rect 565 274248 279575 274648
rect 880 273968 279120 274248
rect 565 273568 279575 273968
rect 880 273288 279120 273568
rect 565 272888 279575 273288
rect 880 272608 279120 272888
rect 565 272208 279575 272608
rect 880 271928 279120 272208
rect 565 271528 279575 271928
rect 880 271248 279120 271528
rect 565 270848 279575 271248
rect 880 270568 279120 270848
rect 565 269488 279575 270568
rect 880 269208 279120 269488
rect 565 268808 279575 269208
rect 880 268528 279120 268808
rect 565 268128 279575 268528
rect 880 267848 279120 268128
rect 565 267448 279575 267848
rect 880 267168 279120 267448
rect 565 266768 279575 267168
rect 880 266488 279120 266768
rect 565 266088 279575 266488
rect 880 265808 279120 266088
rect 565 265408 279575 265808
rect 880 265128 279120 265408
rect 565 264728 279575 265128
rect 880 264448 279120 264728
rect 565 264048 279575 264448
rect 880 263768 279575 264048
rect 565 263368 279575 263768
rect 565 263088 279120 263368
rect 565 262688 279575 263088
rect 880 262408 279120 262688
rect 565 262008 279575 262408
rect 880 261728 279120 262008
rect 565 261328 279575 261728
rect 880 261048 279120 261328
rect 565 260648 279575 261048
rect 880 260368 279120 260648
rect 565 259968 279575 260368
rect 880 259688 279120 259968
rect 565 259288 279575 259688
rect 880 259008 279120 259288
rect 565 258608 279575 259008
rect 880 258328 279120 258608
rect 565 257928 279575 258328
rect 880 257648 279120 257928
rect 565 256568 279575 257648
rect 880 256288 279120 256568
rect 565 255888 279575 256288
rect 880 255608 279120 255888
rect 565 255208 279575 255608
rect 880 254928 279120 255208
rect 565 254528 279575 254928
rect 880 254248 279120 254528
rect 565 253848 279575 254248
rect 880 253568 279120 253848
rect 565 253168 279575 253568
rect 880 252888 279120 253168
rect 565 252488 279575 252888
rect 880 252208 279120 252488
rect 565 251808 279575 252208
rect 880 251528 279120 251808
rect 565 251128 279575 251528
rect 880 250848 279575 251128
rect 565 250448 279575 250848
rect 565 250168 279120 250448
rect 565 249768 279575 250168
rect 880 249488 279120 249768
rect 565 249088 279575 249488
rect 880 248808 279120 249088
rect 565 248408 279575 248808
rect 880 248128 279120 248408
rect 565 247728 279575 248128
rect 880 247448 279120 247728
rect 565 247048 279575 247448
rect 880 246768 279120 247048
rect 565 246368 279575 246768
rect 880 246088 279120 246368
rect 565 245688 279575 246088
rect 880 245408 279120 245688
rect 565 245008 279575 245408
rect 880 244728 279120 245008
rect 565 243648 279575 244728
rect 880 243368 279120 243648
rect 565 242968 279575 243368
rect 880 242688 279120 242968
rect 565 242288 279575 242688
rect 880 242008 279120 242288
rect 565 241608 279575 242008
rect 880 241328 279120 241608
rect 565 240928 279575 241328
rect 880 240648 279120 240928
rect 565 240248 279575 240648
rect 880 239968 279120 240248
rect 565 239568 279575 239968
rect 880 239288 279120 239568
rect 565 238888 279575 239288
rect 880 238608 279120 238888
rect 565 237528 279575 238608
rect 880 237248 279120 237528
rect 565 236848 279575 237248
rect 880 236568 279120 236848
rect 565 236168 279575 236568
rect 880 235888 279120 236168
rect 565 235488 279575 235888
rect 880 235208 279120 235488
rect 565 234808 279575 235208
rect 880 234528 279120 234808
rect 565 234128 279575 234528
rect 880 233848 279120 234128
rect 565 233448 279575 233848
rect 880 233168 279120 233448
rect 565 232768 279575 233168
rect 880 232488 279120 232768
rect 565 232088 279575 232488
rect 880 231808 279120 232088
rect 565 230728 279575 231808
rect 880 230448 279120 230728
rect 565 230048 279575 230448
rect 880 229768 279120 230048
rect 565 229368 279575 229768
rect 880 229088 279120 229368
rect 565 228688 279575 229088
rect 880 228408 279120 228688
rect 565 228008 279575 228408
rect 880 227728 279120 228008
rect 565 227328 279575 227728
rect 880 227048 279120 227328
rect 565 226648 279575 227048
rect 880 226368 279120 226648
rect 565 225968 279575 226368
rect 880 225688 279120 225968
rect 565 224608 279575 225688
rect 880 224328 279120 224608
rect 565 223928 279575 224328
rect 880 223648 279120 223928
rect 565 223248 279575 223648
rect 880 222968 279120 223248
rect 565 222568 279575 222968
rect 880 222288 279120 222568
rect 565 221888 279575 222288
rect 880 221608 279120 221888
rect 565 221208 279575 221608
rect 880 220928 279120 221208
rect 565 220528 279575 220928
rect 880 220248 279120 220528
rect 565 219848 279575 220248
rect 880 219568 279120 219848
rect 565 219168 279575 219568
rect 880 218888 279120 219168
rect 565 217808 279575 218888
rect 880 217528 279120 217808
rect 565 217128 279575 217528
rect 880 216848 279120 217128
rect 565 216448 279575 216848
rect 880 216168 279120 216448
rect 565 215768 279575 216168
rect 880 215488 279120 215768
rect 565 215088 279575 215488
rect 880 214808 279120 215088
rect 565 214408 279575 214808
rect 880 214128 279120 214408
rect 565 213728 279575 214128
rect 880 213448 279120 213728
rect 565 213048 279575 213448
rect 880 212768 279120 213048
rect 565 211688 279575 212768
rect 880 211408 279120 211688
rect 565 211008 279575 211408
rect 880 210728 279120 211008
rect 565 210328 279575 210728
rect 880 210048 279120 210328
rect 565 209648 279575 210048
rect 880 209368 279120 209648
rect 565 208968 279575 209368
rect 880 208688 279120 208968
rect 565 208288 279575 208688
rect 880 208008 279120 208288
rect 565 207608 279575 208008
rect 880 207328 279120 207608
rect 565 206928 279575 207328
rect 880 206648 279120 206928
rect 565 206248 279575 206648
rect 880 205968 279120 206248
rect 565 204888 279575 205968
rect 880 204608 279120 204888
rect 565 204208 279575 204608
rect 880 203928 279120 204208
rect 565 203528 279575 203928
rect 880 203248 279120 203528
rect 565 202848 279575 203248
rect 880 202568 279120 202848
rect 565 202168 279575 202568
rect 880 201888 279120 202168
rect 565 201488 279575 201888
rect 880 201208 279120 201488
rect 565 200808 279575 201208
rect 880 200528 279120 200808
rect 565 200128 279575 200528
rect 880 199848 279120 200128
rect 565 198768 279575 199848
rect 880 198488 279120 198768
rect 565 198088 279575 198488
rect 880 197808 279120 198088
rect 565 197408 279575 197808
rect 880 197128 279120 197408
rect 565 196728 279575 197128
rect 880 196448 279120 196728
rect 565 196048 279575 196448
rect 880 195768 279120 196048
rect 565 195368 279575 195768
rect 880 195088 279120 195368
rect 565 194688 279575 195088
rect 880 194408 279120 194688
rect 565 194008 279575 194408
rect 880 193728 279120 194008
rect 565 193328 279575 193728
rect 880 193048 279575 193328
rect 565 192648 279575 193048
rect 565 192368 279120 192648
rect 565 191968 279575 192368
rect 880 191688 279120 191968
rect 565 191288 279575 191688
rect 880 191008 279120 191288
rect 565 190608 279575 191008
rect 880 190328 279120 190608
rect 565 189928 279575 190328
rect 880 189648 279120 189928
rect 565 189248 279575 189648
rect 880 188968 279120 189248
rect 565 188568 279575 188968
rect 880 188288 279120 188568
rect 565 187888 279575 188288
rect 880 187608 279120 187888
rect 565 187208 279575 187608
rect 880 186928 279120 187208
rect 565 185848 279575 186928
rect 880 185568 279120 185848
rect 565 185168 279575 185568
rect 880 184888 279120 185168
rect 565 184488 279575 184888
rect 880 184208 279120 184488
rect 565 183808 279575 184208
rect 880 183528 279120 183808
rect 565 183128 279575 183528
rect 880 182848 279120 183128
rect 565 182448 279575 182848
rect 880 182168 279120 182448
rect 565 181768 279575 182168
rect 880 181488 279120 181768
rect 565 181088 279575 181488
rect 880 180808 279120 181088
rect 565 180408 279575 180808
rect 880 180128 279575 180408
rect 565 179728 279575 180128
rect 565 179448 279120 179728
rect 565 179048 279575 179448
rect 880 178768 279120 179048
rect 565 178368 279575 178768
rect 880 178088 279120 178368
rect 565 177688 279575 178088
rect 880 177408 279120 177688
rect 565 177008 279575 177408
rect 880 176728 279120 177008
rect 565 176328 279575 176728
rect 880 176048 279120 176328
rect 565 175648 279575 176048
rect 880 175368 279120 175648
rect 565 174968 279575 175368
rect 880 174688 279120 174968
rect 565 174288 279575 174688
rect 880 174008 279120 174288
rect 565 172928 279575 174008
rect 880 172648 279120 172928
rect 565 172248 279575 172648
rect 880 171968 279120 172248
rect 565 171568 279575 171968
rect 880 171288 279120 171568
rect 565 170888 279575 171288
rect 880 170608 279120 170888
rect 565 170208 279575 170608
rect 880 169928 279120 170208
rect 565 169528 279575 169928
rect 880 169248 279120 169528
rect 565 168848 279575 169248
rect 880 168568 279120 168848
rect 565 168168 279575 168568
rect 880 167888 279120 168168
rect 565 167488 279575 167888
rect 880 167208 279575 167488
rect 565 166808 279575 167208
rect 565 166528 279120 166808
rect 565 166128 279575 166528
rect 880 165848 279120 166128
rect 565 165448 279575 165848
rect 880 165168 279120 165448
rect 565 164768 279575 165168
rect 880 164488 279120 164768
rect 565 164088 279575 164488
rect 880 163808 279120 164088
rect 565 163408 279575 163808
rect 880 163128 279120 163408
rect 565 162728 279575 163128
rect 880 162448 279120 162728
rect 565 162048 279575 162448
rect 880 161768 279120 162048
rect 565 161368 279575 161768
rect 880 161088 279120 161368
rect 565 160008 279575 161088
rect 880 159728 279120 160008
rect 565 159328 279575 159728
rect 880 159048 279120 159328
rect 565 158648 279575 159048
rect 880 158368 279120 158648
rect 565 157968 279575 158368
rect 880 157688 279120 157968
rect 565 157288 279575 157688
rect 880 157008 279120 157288
rect 565 156608 279575 157008
rect 880 156328 279120 156608
rect 565 155928 279575 156328
rect 880 155648 279120 155928
rect 565 155248 279575 155648
rect 880 154968 279120 155248
rect 565 153888 279575 154968
rect 880 153608 279120 153888
rect 565 153208 279575 153608
rect 880 152928 279120 153208
rect 565 152528 279575 152928
rect 880 152248 279120 152528
rect 565 151848 279575 152248
rect 880 151568 279120 151848
rect 565 151168 279575 151568
rect 880 150888 279120 151168
rect 565 150488 279575 150888
rect 880 150208 279120 150488
rect 565 149808 279575 150208
rect 880 149528 279120 149808
rect 565 149128 279575 149528
rect 880 148848 279120 149128
rect 565 148448 279575 148848
rect 880 148168 279120 148448
rect 565 147088 279575 148168
rect 880 146808 279120 147088
rect 565 146408 279575 146808
rect 880 146128 279120 146408
rect 565 145728 279575 146128
rect 880 145448 279120 145728
rect 565 145048 279575 145448
rect 880 144768 279120 145048
rect 565 144368 279575 144768
rect 880 144088 279120 144368
rect 565 143688 279575 144088
rect 880 143408 279120 143688
rect 565 143008 279575 143408
rect 880 142728 279120 143008
rect 565 142328 279575 142728
rect 880 142048 279120 142328
rect 565 140968 279575 142048
rect 880 140688 279120 140968
rect 565 140288 279575 140688
rect 880 140008 279120 140288
rect 565 139608 279575 140008
rect 880 139328 279120 139608
rect 565 138928 279575 139328
rect 880 138648 279120 138928
rect 565 138248 279575 138648
rect 880 137968 279120 138248
rect 565 137568 279575 137968
rect 880 137288 279120 137568
rect 565 136888 279575 137288
rect 880 136608 279120 136888
rect 565 136208 279575 136608
rect 880 135928 279120 136208
rect 565 135528 279575 135928
rect 880 135248 279120 135528
rect 565 134168 279575 135248
rect 880 133888 279120 134168
rect 565 133488 279575 133888
rect 880 133208 279120 133488
rect 565 132808 279575 133208
rect 880 132528 279120 132808
rect 565 132128 279575 132528
rect 880 131848 279120 132128
rect 565 131448 279575 131848
rect 880 131168 279120 131448
rect 565 130768 279575 131168
rect 880 130488 279120 130768
rect 565 130088 279575 130488
rect 880 129808 279120 130088
rect 565 129408 279575 129808
rect 880 129128 279120 129408
rect 565 128048 279575 129128
rect 880 127768 279120 128048
rect 565 127368 279575 127768
rect 880 127088 279120 127368
rect 565 126688 279575 127088
rect 880 126408 279120 126688
rect 565 126008 279575 126408
rect 880 125728 279120 126008
rect 565 125328 279575 125728
rect 880 125048 279120 125328
rect 565 124648 279575 125048
rect 880 124368 279120 124648
rect 565 123968 279575 124368
rect 880 123688 279120 123968
rect 565 123288 279575 123688
rect 880 123008 279120 123288
rect 565 122608 279575 123008
rect 880 122328 279120 122608
rect 565 121248 279575 122328
rect 880 120968 279120 121248
rect 565 120568 279575 120968
rect 880 120288 279120 120568
rect 565 119888 279575 120288
rect 880 119608 279120 119888
rect 565 119208 279575 119608
rect 880 118928 279120 119208
rect 565 118528 279575 118928
rect 880 118248 279120 118528
rect 565 117848 279575 118248
rect 880 117568 279120 117848
rect 565 117168 279575 117568
rect 880 116888 279120 117168
rect 565 116488 279575 116888
rect 880 116208 279120 116488
rect 565 115128 279575 116208
rect 880 114848 279120 115128
rect 565 114448 279575 114848
rect 880 114168 279120 114448
rect 565 113768 279575 114168
rect 880 113488 279120 113768
rect 565 113088 279575 113488
rect 880 112808 279120 113088
rect 565 112408 279575 112808
rect 880 112128 279120 112408
rect 565 111728 279575 112128
rect 880 111448 279120 111728
rect 565 111048 279575 111448
rect 880 110768 279120 111048
rect 565 110368 279575 110768
rect 880 110088 279120 110368
rect 565 109688 279575 110088
rect 880 109408 279575 109688
rect 565 109008 279575 109408
rect 565 108728 279120 109008
rect 565 108328 279575 108728
rect 880 108048 279120 108328
rect 565 107648 279575 108048
rect 880 107368 279120 107648
rect 565 106968 279575 107368
rect 880 106688 279120 106968
rect 565 106288 279575 106688
rect 880 106008 279120 106288
rect 565 105608 279575 106008
rect 880 105328 279120 105608
rect 565 104928 279575 105328
rect 880 104648 279120 104928
rect 565 104248 279575 104648
rect 880 103968 279120 104248
rect 565 103568 279575 103968
rect 880 103288 279120 103568
rect 565 102208 279575 103288
rect 880 101928 279120 102208
rect 565 101528 279575 101928
rect 880 101248 279120 101528
rect 565 100848 279575 101248
rect 880 100568 279120 100848
rect 565 100168 279575 100568
rect 880 99888 279120 100168
rect 565 99488 279575 99888
rect 880 99208 279120 99488
rect 565 98808 279575 99208
rect 880 98528 279120 98808
rect 565 98128 279575 98528
rect 880 97848 279120 98128
rect 565 97448 279575 97848
rect 880 97168 279120 97448
rect 565 96768 279575 97168
rect 880 96488 279575 96768
rect 565 96088 279575 96488
rect 565 95808 279120 96088
rect 565 95408 279575 95808
rect 880 95128 279120 95408
rect 565 94728 279575 95128
rect 880 94448 279120 94728
rect 565 94048 279575 94448
rect 880 93768 279120 94048
rect 565 93368 279575 93768
rect 880 93088 279120 93368
rect 565 92688 279575 93088
rect 880 92408 279120 92688
rect 565 92008 279575 92408
rect 880 91728 279120 92008
rect 565 91328 279575 91728
rect 880 91048 279120 91328
rect 565 90648 279575 91048
rect 880 90368 279120 90648
rect 565 89288 279575 90368
rect 880 89008 279120 89288
rect 565 88608 279575 89008
rect 880 88328 279120 88608
rect 565 87928 279575 88328
rect 880 87648 279120 87928
rect 565 87248 279575 87648
rect 880 86968 279120 87248
rect 565 86568 279575 86968
rect 880 86288 279120 86568
rect 565 85888 279575 86288
rect 880 85608 279120 85888
rect 565 85208 279575 85608
rect 880 84928 279120 85208
rect 565 84528 279575 84928
rect 880 84248 279120 84528
rect 565 83848 279575 84248
rect 880 83568 279575 83848
rect 565 83168 279575 83568
rect 565 82888 279120 83168
rect 565 82488 279575 82888
rect 880 82208 279120 82488
rect 565 81808 279575 82208
rect 880 81528 279120 81808
rect 565 81128 279575 81528
rect 880 80848 279120 81128
rect 565 80448 279575 80848
rect 880 80168 279120 80448
rect 565 79768 279575 80168
rect 880 79488 279120 79768
rect 565 79088 279575 79488
rect 880 78808 279120 79088
rect 565 78408 279575 78808
rect 880 78128 279120 78408
rect 565 77728 279575 78128
rect 880 77448 279120 77728
rect 565 76368 279575 77448
rect 880 76088 279120 76368
rect 565 75688 279575 76088
rect 880 75408 279120 75688
rect 565 75008 279575 75408
rect 880 74728 279120 75008
rect 565 74328 279575 74728
rect 880 74048 279120 74328
rect 565 73648 279575 74048
rect 880 73368 279120 73648
rect 565 72968 279575 73368
rect 880 72688 279120 72968
rect 565 72288 279575 72688
rect 880 72008 279120 72288
rect 565 71608 279575 72008
rect 880 71328 279120 71608
rect 565 70248 279575 71328
rect 880 69968 279120 70248
rect 565 69568 279575 69968
rect 880 69288 279120 69568
rect 565 68888 279575 69288
rect 880 68608 279120 68888
rect 565 68208 279575 68608
rect 880 67928 279120 68208
rect 565 67528 279575 67928
rect 880 67248 279120 67528
rect 565 66848 279575 67248
rect 880 66568 279120 66848
rect 565 66168 279575 66568
rect 880 65888 279120 66168
rect 565 65488 279575 65888
rect 880 65208 279120 65488
rect 565 64808 279575 65208
rect 880 64528 279120 64808
rect 565 63448 279575 64528
rect 880 63168 279120 63448
rect 565 62768 279575 63168
rect 880 62488 279120 62768
rect 565 62088 279575 62488
rect 880 61808 279120 62088
rect 565 61408 279575 61808
rect 880 61128 279120 61408
rect 565 60728 279575 61128
rect 880 60448 279120 60728
rect 565 60048 279575 60448
rect 880 59768 279120 60048
rect 565 59368 279575 59768
rect 880 59088 279120 59368
rect 565 58688 279575 59088
rect 880 58408 279120 58688
rect 565 57328 279575 58408
rect 880 57048 279120 57328
rect 565 56648 279575 57048
rect 880 56368 279120 56648
rect 565 55968 279575 56368
rect 880 55688 279120 55968
rect 565 55288 279575 55688
rect 880 55008 279120 55288
rect 565 54608 279575 55008
rect 880 54328 279120 54608
rect 565 53928 279575 54328
rect 880 53648 279120 53928
rect 565 53248 279575 53648
rect 880 52968 279120 53248
rect 565 52568 279575 52968
rect 880 52288 279120 52568
rect 565 51888 279575 52288
rect 880 51608 279120 51888
rect 565 50528 279575 51608
rect 880 50248 279120 50528
rect 565 49848 279575 50248
rect 880 49568 279120 49848
rect 565 49168 279575 49568
rect 880 48888 279120 49168
rect 565 48488 279575 48888
rect 880 48208 279120 48488
rect 565 47808 279575 48208
rect 880 47528 279120 47808
rect 565 47128 279575 47528
rect 880 46848 279120 47128
rect 565 46448 279575 46848
rect 880 46168 279120 46448
rect 565 45768 279575 46168
rect 880 45488 279120 45768
rect 565 44408 279575 45488
rect 880 44128 279120 44408
rect 565 43728 279575 44128
rect 880 43448 279120 43728
rect 565 43048 279575 43448
rect 880 42768 279120 43048
rect 565 42368 279575 42768
rect 880 42088 279120 42368
rect 565 41688 279575 42088
rect 880 41408 279120 41688
rect 565 41008 279575 41408
rect 880 40728 279120 41008
rect 565 40328 279575 40728
rect 880 40048 279120 40328
rect 565 39648 279575 40048
rect 880 39368 279120 39648
rect 565 38968 279575 39368
rect 880 38688 279120 38968
rect 565 37608 279575 38688
rect 880 37328 279120 37608
rect 565 36928 279575 37328
rect 880 36648 279120 36928
rect 565 36248 279575 36648
rect 880 35968 279120 36248
rect 565 35568 279575 35968
rect 880 35288 279120 35568
rect 565 34888 279575 35288
rect 880 34608 279120 34888
rect 565 34208 279575 34608
rect 880 33928 279120 34208
rect 565 33528 279575 33928
rect 880 33248 279120 33528
rect 565 32848 279575 33248
rect 880 32568 279120 32848
rect 565 31488 279575 32568
rect 880 31208 279120 31488
rect 565 30808 279575 31208
rect 880 30528 279120 30808
rect 565 30128 279575 30528
rect 880 29848 279120 30128
rect 565 29448 279575 29848
rect 880 29168 279120 29448
rect 565 28768 279575 29168
rect 880 28488 279120 28768
rect 565 28088 279575 28488
rect 880 27808 279120 28088
rect 565 27408 279575 27808
rect 880 27128 279120 27408
rect 565 26728 279575 27128
rect 880 26448 279120 26728
rect 565 26048 279575 26448
rect 880 25768 279575 26048
rect 565 25368 279575 25768
rect 565 25088 279120 25368
rect 565 24688 279575 25088
rect 880 24408 279120 24688
rect 565 24008 279575 24408
rect 880 23728 279120 24008
rect 565 23328 279575 23728
rect 880 23048 279120 23328
rect 565 22648 279575 23048
rect 880 22368 279120 22648
rect 565 21968 279575 22368
rect 880 21688 279120 21968
rect 565 21288 279575 21688
rect 880 21008 279120 21288
rect 565 20608 279575 21008
rect 880 20328 279120 20608
rect 565 19928 279575 20328
rect 880 19648 279120 19928
rect 565 18568 279575 19648
rect 880 18288 279120 18568
rect 565 17888 279575 18288
rect 880 17608 279120 17888
rect 565 17208 279575 17608
rect 880 16928 279120 17208
rect 565 16528 279575 16928
rect 880 16248 279120 16528
rect 565 15848 279575 16248
rect 880 15568 279120 15848
rect 565 15168 279575 15568
rect 880 14888 279120 15168
rect 565 14488 279575 14888
rect 880 14208 279120 14488
rect 565 13808 279575 14208
rect 880 13528 279120 13808
rect 565 13128 279575 13528
rect 880 12848 279575 13128
rect 565 12448 279575 12848
rect 565 12168 279120 12448
rect 565 11768 279575 12168
rect 880 11488 279120 11768
rect 565 11088 279575 11488
rect 880 10808 279120 11088
rect 565 10408 279575 10808
rect 880 10128 279120 10408
rect 565 9728 279575 10128
rect 880 9448 279120 9728
rect 565 9048 279575 9448
rect 880 8768 279120 9048
rect 565 8368 279575 8768
rect 880 8088 279120 8368
rect 565 7688 279575 8088
rect 880 7408 279120 7688
rect 565 7008 279575 7408
rect 880 6728 279120 7008
rect 565 5648 279575 6728
rect 880 5368 279120 5648
rect 565 4968 279575 5368
rect 880 4688 279120 4968
rect 565 4288 279575 4688
rect 880 4008 279120 4288
rect 565 3608 279575 4008
rect 880 3328 279120 3608
rect 565 2928 279575 3328
rect 880 2648 279120 2928
rect 565 2248 279575 2648
rect 880 1968 279120 2248
rect 565 1568 279575 1968
rect 880 1288 279120 1568
rect 565 888 279575 1288
rect 880 715 279120 888
<< metal4 >>
rect 4208 2128 4528 357456
rect 19568 2128 19888 357456
rect 34928 2128 35248 357456
rect 50288 2128 50608 357456
rect 65648 2128 65968 357456
rect 81008 2128 81328 357456
rect 96368 2128 96688 357456
rect 111728 2128 112048 357456
rect 127088 2128 127408 357456
rect 142448 2128 142768 357456
rect 157808 2128 158128 357456
rect 173168 2128 173488 357456
rect 188528 2128 188848 357456
rect 203888 2128 204208 357456
rect 219248 2128 219568 357456
rect 234608 2128 234928 357456
rect 249968 2128 250288 357456
rect 265328 2128 265648 357456
<< obsm4 >>
rect 611 2048 4128 357237
rect 4608 2048 19488 357237
rect 19968 2048 34848 357237
rect 35328 2048 50208 357237
rect 50688 2048 65568 357237
rect 66048 2048 80928 357237
rect 81408 2048 96288 357237
rect 96768 2048 111648 357237
rect 112128 2048 127008 357237
rect 127488 2048 142368 357237
rect 142848 2048 157728 357237
rect 158208 2048 173088 357237
rect 173568 2048 188448 357237
rect 188928 2048 203808 357237
rect 204288 2048 219168 357237
rect 219648 2048 234528 357237
rect 235008 2048 249888 357237
rect 250368 2048 265248 357237
rect 265728 2048 277229 357237
rect 611 1531 277229 2048
<< labels >>
rlabel metal3 s 279200 23128 280000 23248 6 boot_addr_i[0]
port 1 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 boot_addr_i[10]
port 2 nsew signal input
rlabel metal3 s 0 212848 800 212968 6 boot_addr_i[11]
port 3 nsew signal input
rlabel metal3 s 0 331168 800 331288 6 boot_addr_i[12]
port 4 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 boot_addr_i[13]
port 5 nsew signal input
rlabel metal2 s 278226 0 278282 800 6 boot_addr_i[14]
port 6 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 boot_addr_i[15]
port 7 nsew signal input
rlabel metal3 s 0 220328 800 220448 6 boot_addr_i[16]
port 8 nsew signal input
rlabel metal3 s 279200 87048 280000 87168 6 boot_addr_i[17]
port 9 nsew signal input
rlabel metal3 s 0 337288 800 337408 6 boot_addr_i[18]
port 10 nsew signal input
rlabel metal3 s 0 189048 800 189168 6 boot_addr_i[19]
port 11 nsew signal input
rlabel metal3 s 0 278128 800 278248 6 boot_addr_i[1]
port 12 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 boot_addr_i[20]
port 13 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 boot_addr_i[21]
port 14 nsew signal input
rlabel metal3 s 279200 307368 280000 307488 6 boot_addr_i[22]
port 15 nsew signal input
rlabel metal2 s 17406 359200 17462 360000 6 boot_addr_i[23]
port 16 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 boot_addr_i[24]
port 17 nsew signal input
rlabel metal3 s 279200 10208 280000 10328 6 boot_addr_i[25]
port 18 nsew signal input
rlabel metal2 s 14830 359200 14886 360000 6 boot_addr_i[26]
port 19 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 boot_addr_i[27]
port 20 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 boot_addr_i[28]
port 21 nsew signal input
rlabel metal2 s 39302 359200 39358 360000 6 boot_addr_i[29]
port 22 nsew signal input
rlabel metal3 s 0 168648 800 168768 6 boot_addr_i[2]
port 23 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 boot_addr_i[30]
port 24 nsew signal input
rlabel metal3 s 0 248888 800 249008 6 boot_addr_i[31]
port 25 nsew signal input
rlabel metal2 s 207386 0 207442 800 6 boot_addr_i[3]
port 26 nsew signal input
rlabel metal3 s 279200 1368 280000 1488 6 boot_addr_i[4]
port 27 nsew signal input
rlabel metal3 s 0 290368 800 290488 6 boot_addr_i[5]
port 28 nsew signal input
rlabel metal3 s 279200 114248 280000 114368 6 boot_addr_i[6]
port 29 nsew signal input
rlabel metal3 s 279200 197208 280000 197328 6 boot_addr_i[7]
port 30 nsew signal input
rlabel metal3 s 279200 27208 280000 27328 6 boot_addr_i[8]
port 31 nsew signal input
rlabel metal3 s 279200 269288 280000 269408 6 boot_addr_i[9]
port 32 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 clk
port 33 nsew signal input
rlabel metal2 s 185490 359200 185546 360000 6 clock_gating_i
port 34 nsew signal input
rlabel metal3 s 279200 46248 280000 46368 6 core_busy_o
port 35 nsew signal output
rlabel metal2 s 130106 359200 130162 360000 6 core_master_ar_addr[0]
port 36 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 core_master_ar_addr[10]
port 37 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 core_master_ar_addr[11]
port 38 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 core_master_ar_addr[12]
port 39 nsew signal output
rlabel metal2 s 196438 0 196494 800 6 core_master_ar_addr[13]
port 40 nsew signal output
rlabel metal3 s 0 328448 800 328568 6 core_master_ar_addr[14]
port 41 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 core_master_ar_addr[15]
port 42 nsew signal output
rlabel metal2 s 229926 0 229982 800 6 core_master_ar_addr[16]
port 43 nsew signal output
rlabel metal3 s 0 347488 800 347608 6 core_master_ar_addr[17]
port 44 nsew signal output
rlabel metal3 s 279200 256368 280000 256488 6 core_master_ar_addr[18]
port 45 nsew signal output
rlabel metal2 s 104346 359200 104402 360000 6 core_master_ar_addr[19]
port 46 nsew signal output
rlabel metal3 s 0 251608 800 251728 6 core_master_ar_addr[1]
port 47 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 core_master_ar_addr[20]
port 48 nsew signal output
rlabel metal3 s 279200 120368 280000 120488 6 core_master_ar_addr[21]
port 49 nsew signal output
rlabel metal3 s 279200 291048 280000 291168 6 core_master_ar_addr[22]
port 50 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 core_master_ar_addr[23]
port 51 nsew signal output
rlabel metal2 s 241518 359200 241574 360000 6 core_master_ar_addr[24]
port 52 nsew signal output
rlabel metal2 s 232502 0 232558 800 6 core_master_ar_addr[25]
port 53 nsew signal output
rlabel metal3 s 279200 303968 280000 304088 6 core_master_ar_addr[26]
port 54 nsew signal output
rlabel metal3 s 0 343408 800 343528 6 core_master_ar_addr[27]
port 55 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 core_master_ar_addr[28]
port 56 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 core_master_ar_addr[29]
port 57 nsew signal output
rlabel metal2 s 56046 359200 56102 360000 6 core_master_ar_addr[2]
port 58 nsew signal output
rlabel metal3 s 279200 45568 280000 45688 6 core_master_ar_addr[30]
port 59 nsew signal output
rlabel metal3 s 0 195168 800 195288 6 core_master_ar_addr[31]
port 60 nsew signal output
rlabel metal3 s 279200 145528 280000 145648 6 core_master_ar_addr[3]
port 61 nsew signal output
rlabel metal3 s 279200 286288 280000 286408 6 core_master_ar_addr[4]
port 62 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 core_master_ar_addr[5]
port 63 nsew signal output
rlabel metal3 s 279200 182248 280000 182368 6 core_master_ar_addr[6]
port 64 nsew signal output
rlabel metal3 s 0 329808 800 329928 6 core_master_ar_addr[7]
port 65 nsew signal output
rlabel metal2 s 233146 0 233202 800 6 core_master_ar_addr[8]
port 66 nsew signal output
rlabel metal2 s 72146 359200 72202 360000 6 core_master_ar_addr[9]
port 67 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 core_master_ar_burst[0]
port 68 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 core_master_ar_burst[1]
port 69 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 core_master_ar_cache[0]
port 70 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 core_master_ar_cache[1]
port 71 nsew signal output
rlabel metal3 s 0 270648 800 270768 6 core_master_ar_cache[2]
port 72 nsew signal output
rlabel metal3 s 279200 295128 280000 295248 6 core_master_ar_cache[3]
port 73 nsew signal output
rlabel metal3 s 279200 274728 280000 274848 6 core_master_ar_id[0]
port 74 nsew signal output
rlabel metal3 s 0 348848 800 348968 6 core_master_ar_id[1]
port 75 nsew signal output
rlabel metal3 s 279200 210808 280000 210928 6 core_master_ar_id[2]
port 76 nsew signal output
rlabel metal2 s 150070 359200 150126 360000 6 core_master_ar_id[3]
port 77 nsew signal output
rlabel metal3 s 279200 8168 280000 8288 6 core_master_ar_id[4]
port 78 nsew signal output
rlabel metal3 s 0 142128 800 142248 6 core_master_ar_id[5]
port 79 nsew signal output
rlabel metal3 s 279200 62568 280000 62688 6 core_master_ar_id[6]
port 80 nsew signal output
rlabel metal2 s 186778 359200 186834 360000 6 core_master_ar_id[7]
port 81 nsew signal output
rlabel metal3 s 0 280848 800 280968 6 core_master_ar_id[8]
port 82 nsew signal output
rlabel metal2 s 62486 359200 62542 360000 6 core_master_ar_id[9]
port 83 nsew signal output
rlabel metal2 s 142342 359200 142398 360000 6 core_master_ar_len[0]
port 84 nsew signal output
rlabel metal3 s 0 297848 800 297968 6 core_master_ar_len[1]
port 85 nsew signal output
rlabel metal3 s 279200 16328 280000 16448 6 core_master_ar_len[2]
port 86 nsew signal output
rlabel metal2 s 24490 359200 24546 360000 6 core_master_ar_len[3]
port 87 nsew signal output
rlabel metal2 s 256974 0 257030 800 6 core_master_ar_len[4]
port 88 nsew signal output
rlabel metal3 s 279200 204008 280000 204128 6 core_master_ar_len[5]
port 89 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 core_master_ar_len[6]
port 90 nsew signal output
rlabel metal2 s 35438 359200 35494 360000 6 core_master_ar_len[7]
port 91 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 core_master_ar_lock
port 92 nsew signal output
rlabel metal3 s 279200 259768 280000 259888 6 core_master_ar_prot[0]
port 93 nsew signal output
rlabel metal2 s 199014 0 199070 800 6 core_master_ar_prot[1]
port 94 nsew signal output
rlabel metal2 s 184846 359200 184902 360000 6 core_master_ar_prot[2]
port 95 nsew signal output
rlabel metal2 s 25778 359200 25834 360000 6 core_master_ar_qos[0]
port 96 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 core_master_ar_qos[1]
port 97 nsew signal output
rlabel metal3 s 279200 136688 280000 136808 6 core_master_ar_qos[2]
port 98 nsew signal output
rlabel metal2 s 64418 359200 64474 360000 6 core_master_ar_qos[3]
port 99 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 core_master_ar_ready
port 100 nsew signal input
rlabel metal3 s 279200 127168 280000 127288 6 core_master_ar_region[0]
port 101 nsew signal output
rlabel metal2 s 202878 359200 202934 360000 6 core_master_ar_region[1]
port 102 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 core_master_ar_region[2]
port 103 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 core_master_ar_region[3]
port 104 nsew signal output
rlabel metal3 s 279200 293088 280000 293208 6 core_master_ar_size[0]
port 105 nsew signal output
rlabel metal3 s 0 287648 800 287768 6 core_master_ar_size[1]
port 106 nsew signal output
rlabel metal3 s 279200 221008 280000 221128 6 core_master_ar_size[2]
port 107 nsew signal output
rlabel metal3 s 0 180888 800 181008 6 core_master_ar_user[-1]
port 108 nsew signal output
rlabel metal3 s 279200 352928 280000 353048 6 core_master_ar_user[0]
port 109 nsew signal output
rlabel metal3 s 0 219648 800 219768 6 core_master_ar_valid
port 110 nsew signal output
rlabel metal3 s 0 244808 800 244928 6 core_master_aw_addr[0]
port 111 nsew signal output
rlabel metal3 s 279200 131928 280000 132048 6 core_master_aw_addr[10]
port 112 nsew signal output
rlabel metal3 s 0 333208 800 333328 6 core_master_aw_addr[11]
port 113 nsew signal output
rlabel metal3 s 279200 223728 280000 223848 6 core_master_aw_addr[12]
port 114 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 core_master_aw_addr[13]
port 115 nsew signal output
rlabel metal2 s 264702 359200 264758 360000 6 core_master_aw_addr[14]
port 116 nsew signal output
rlabel metal3 s 279200 213528 280000 213648 6 core_master_aw_addr[15]
port 117 nsew signal output
rlabel metal3 s 279200 261128 280000 261248 6 core_master_aw_addr[16]
port 118 nsew signal output
rlabel metal3 s 279200 42168 280000 42288 6 core_master_aw_addr[17]
port 119 nsew signal output
rlabel metal2 s 222198 359200 222254 360000 6 core_master_aw_addr[18]
port 120 nsew signal output
rlabel metal3 s 279200 318928 280000 319048 6 core_master_aw_addr[19]
port 121 nsew signal output
rlabel metal2 s 124954 359200 125010 360000 6 core_master_aw_addr[1]
port 122 nsew signal output
rlabel metal2 s 230570 359200 230626 360000 6 core_master_aw_addr[20]
port 123 nsew signal output
rlabel metal3 s 279200 335248 280000 335368 6 core_master_aw_addr[21]
port 124 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 core_master_aw_addr[22]
port 125 nsew signal output
rlabel metal3 s 279200 30608 280000 30728 6 core_master_aw_addr[23]
port 126 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 core_master_aw_addr[24]
port 127 nsew signal output
rlabel metal2 s 258906 359200 258962 360000 6 core_master_aw_addr[25]
port 128 nsew signal output
rlabel metal3 s 279200 22448 280000 22568 6 core_master_aw_addr[26]
port 129 nsew signal output
rlabel metal3 s 0 182928 800 183048 6 core_master_aw_addr[27]
port 130 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 core_master_aw_addr[28]
port 131 nsew signal output
rlabel metal2 s 170678 359200 170734 360000 6 core_master_aw_addr[29]
port 132 nsew signal output
rlabel metal2 s 253754 359200 253810 360000 6 core_master_aw_addr[2]
port 133 nsew signal output
rlabel metal3 s 279200 220328 280000 220448 6 core_master_aw_addr[30]
port 134 nsew signal output
rlabel metal2 s 266634 359200 266690 360000 6 core_master_aw_addr[31]
port 135 nsew signal output
rlabel metal3 s 279200 73448 280000 73568 6 core_master_aw_addr[3]
port 136 nsew signal output
rlabel metal2 s 167458 359200 167514 360000 6 core_master_aw_addr[4]
port 137 nsew signal output
rlabel metal3 s 279200 2048 280000 2168 6 core_master_aw_addr[5]
port 138 nsew signal output
rlabel metal2 s 218334 0 218390 800 6 core_master_aw_addr[6]
port 139 nsew signal output
rlabel metal3 s 279200 230528 280000 230648 6 core_master_aw_addr[7]
port 140 nsew signal output
rlabel metal2 s 231858 359200 231914 360000 6 core_master_aw_addr[8]
port 141 nsew signal output
rlabel metal2 s 264702 0 264758 800 6 core_master_aw_addr[9]
port 142 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 core_master_aw_burst[0]
port 143 nsew signal output
rlabel metal3 s 279200 210128 280000 210248 6 core_master_aw_burst[1]
port 144 nsew signal output
rlabel metal3 s 279200 349528 280000 349648 6 core_master_aw_cache[0]
port 145 nsew signal output
rlabel metal2 s 202234 359200 202290 360000 6 core_master_aw_cache[1]
port 146 nsew signal output
rlabel metal2 s 65706 359200 65762 360000 6 core_master_aw_cache[2]
port 147 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 core_master_aw_cache[3]
port 148 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 core_master_aw_id[0]
port 149 nsew signal output
rlabel metal3 s 279200 59848 280000 59968 6 core_master_aw_id[1]
port 150 nsew signal output
rlabel metal3 s 279200 325728 280000 325848 6 core_master_aw_id[2]
port 151 nsew signal output
rlabel metal3 s 0 312808 800 312928 6 core_master_aw_id[3]
port 152 nsew signal output
rlabel metal3 s 279200 315528 280000 315648 6 core_master_aw_id[4]
port 153 nsew signal output
rlabel metal3 s 279200 342728 280000 342848 6 core_master_aw_id[5]
port 154 nsew signal output
rlabel metal3 s 0 208088 800 208208 6 core_master_aw_id[6]
port 155 nsew signal output
rlabel metal3 s 0 314168 800 314288 6 core_master_aw_id[7]
port 156 nsew signal output
rlabel metal3 s 279200 110848 280000 110968 6 core_master_aw_id[8]
port 157 nsew signal output
rlabel metal2 s 262126 0 262182 800 6 core_master_aw_id[9]
port 158 nsew signal output
rlabel metal3 s 279200 185648 280000 185768 6 core_master_aw_len[0]
port 159 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 core_master_aw_len[1]
port 160 nsew signal output
rlabel metal2 s 239586 0 239642 800 6 core_master_aw_len[2]
port 161 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 core_master_aw_len[3]
port 162 nsew signal output
rlabel metal3 s 0 247528 800 247648 6 core_master_aw_len[4]
port 163 nsew signal output
rlabel metal3 s 279200 302608 280000 302728 6 core_master_aw_len[5]
port 164 nsew signal output
rlabel metal3 s 0 323688 800 323808 6 core_master_aw_len[6]
port 165 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 core_master_aw_len[7]
port 166 nsew signal output
rlabel metal3 s 0 193808 800 193928 6 core_master_aw_lock
port 167 nsew signal output
rlabel metal2 s 202878 0 202934 800 6 core_master_aw_prot[0]
port 168 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 core_master_aw_prot[1]
port 169 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 core_master_aw_prot[2]
port 170 nsew signal output
rlabel metal3 s 279200 85688 280000 85808 6 core_master_aw_qos[0]
port 171 nsew signal output
rlabel metal3 s 0 323008 800 323128 6 core_master_aw_qos[1]
port 172 nsew signal output
rlabel metal3 s 279200 129208 280000 129328 6 core_master_aw_qos[2]
port 173 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 core_master_aw_qos[3]
port 174 nsew signal output
rlabel metal3 s 0 288328 800 288448 6 core_master_aw_ready
port 175 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 core_master_aw_region[0]
port 176 nsew signal output
rlabel metal2 s 131394 359200 131450 360000 6 core_master_aw_region[1]
port 177 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 core_master_aw_region[2]
port 178 nsew signal output
rlabel metal2 s 21270 359200 21326 360000 6 core_master_aw_region[3]
port 179 nsew signal output
rlabel metal3 s 279200 116968 280000 117088 6 core_master_aw_size[0]
port 180 nsew signal output
rlabel metal3 s 279200 267928 280000 268048 6 core_master_aw_size[1]
port 181 nsew signal output
rlabel metal3 s 279200 254328 280000 254448 6 core_master_aw_size[2]
port 182 nsew signal output
rlabel metal3 s 279200 119688 280000 119808 6 core_master_aw_user[-1]
port 183 nsew signal output
rlabel metal3 s 279200 165248 280000 165368 6 core_master_aw_user[0]
port 184 nsew signal output
rlabel metal3 s 279200 121048 280000 121168 6 core_master_aw_valid
port 185 nsew signal output
rlabel metal2 s 227994 0 228050 800 6 core_master_b_id[0]
port 186 nsew signal input
rlabel metal2 s 102414 359200 102470 360000 6 core_master_b_id[1]
port 187 nsew signal input
rlabel metal2 s 169390 359200 169446 360000 6 core_master_b_id[2]
port 188 nsew signal input
rlabel metal2 s 53470 359200 53526 360000 6 core_master_b_id[3]
port 189 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 core_master_b_id[4]
port 190 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 core_master_b_id[5]
port 191 nsew signal input
rlabel metal2 s 20626 359200 20682 360000 6 core_master_b_id[6]
port 192 nsew signal input
rlabel metal2 s 99194 359200 99250 360000 6 core_master_b_id[7]
port 193 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 core_master_b_id[8]
port 194 nsew signal input
rlabel metal3 s 279200 229848 280000 229968 6 core_master_b_id[9]
port 195 nsew signal input
rlabel metal3 s 279200 166608 280000 166728 6 core_master_b_ready
port 196 nsew signal output
rlabel metal3 s 0 227128 800 227248 6 core_master_b_resp[0]
port 197 nsew signal input
rlabel metal3 s 279200 155728 280000 155848 6 core_master_b_resp[1]
port 198 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 core_master_b_user[-1]
port 199 nsew signal input
rlabel metal2 s 192574 359200 192630 360000 6 core_master_b_user[0]
port 200 nsew signal input
rlabel metal3 s 279200 252288 280000 252408 6 core_master_b_valid
port 201 nsew signal input
rlabel metal2 s 173254 359200 173310 360000 6 core_master_r_data[0]
port 202 nsew signal input
rlabel metal2 s 124310 359200 124366 360000 6 core_master_r_data[10]
port 203 nsew signal input
rlabel metal3 s 0 190408 800 190528 6 core_master_r_data[11]
port 204 nsew signal input
rlabel metal2 s 95974 359200 96030 360000 6 core_master_r_data[12]
port 205 nsew signal input
rlabel metal3 s 0 229168 800 229288 6 core_master_r_data[13]
port 206 nsew signal input
rlabel metal3 s 0 352248 800 352368 6 core_master_r_data[14]
port 207 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 core_master_r_data[15]
port 208 nsew signal input
rlabel metal3 s 0 221688 800 221808 6 core_master_r_data[16]
port 209 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 core_master_r_data[17]
port 210 nsew signal input
rlabel metal2 s 174542 359200 174598 360000 6 core_master_r_data[18]
port 211 nsew signal input
rlabel metal2 s 275650 0 275706 800 6 core_master_r_data[19]
port 212 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 core_master_r_data[1]
port 213 nsew signal input
rlabel metal3 s 0 265888 800 266008 6 core_master_r_data[20]
port 214 nsew signal input
rlabel metal3 s 0 272688 800 272808 6 core_master_r_data[21]
port 215 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 core_master_r_data[22]
port 216 nsew signal input
rlabel metal2 s 249890 359200 249946 360000 6 core_master_r_data[23]
port 217 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 core_master_r_data[24]
port 218 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 core_master_r_data[25]
port 219 nsew signal input
rlabel metal2 s 94686 359200 94742 360000 6 core_master_r_data[26]
port 220 nsew signal input
rlabel metal3 s 279200 48968 280000 49088 6 core_master_r_data[27]
port 221 nsew signal input
rlabel metal3 s 279200 17008 280000 17128 6 core_master_r_data[28]
port 222 nsew signal input
rlabel metal2 s 256330 359200 256386 360000 6 core_master_r_data[29]
port 223 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 core_master_r_data[2]
port 224 nsew signal input
rlabel metal3 s 279200 116288 280000 116408 6 core_master_r_data[30]
port 225 nsew signal input
rlabel metal3 s 0 200608 800 200728 6 core_master_r_data[31]
port 226 nsew signal input
rlabel metal3 s 279200 165928 280000 166048 6 core_master_r_data[32]
port 227 nsew signal input
rlabel metal2 s 183558 359200 183614 360000 6 core_master_r_data[33]
port 228 nsew signal input
rlabel metal2 s 26422 359200 26478 360000 6 core_master_r_data[34]
port 229 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 core_master_r_data[35]
port 230 nsew signal input
rlabel metal2 s 161018 359200 161074 360000 6 core_master_r_data[36]
port 231 nsew signal input
rlabel metal3 s 0 234608 800 234728 6 core_master_r_data[37]
port 232 nsew signal input
rlabel metal3 s 279200 163208 280000 163328 6 core_master_r_data[38]
port 233 nsew signal input
rlabel metal2 s 40590 359200 40646 360000 6 core_master_r_data[39]
port 234 nsew signal input
rlabel metal3 s 279200 177488 280000 177608 6 core_master_r_data[3]
port 235 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 core_master_r_data[40]
port 236 nsew signal input
rlabel metal3 s 279200 139408 280000 139528 6 core_master_r_data[41]
port 237 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 core_master_r_data[42]
port 238 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 core_master_r_data[43]
port 239 nsew signal input
rlabel metal2 s 222842 359200 222898 360000 6 core_master_r_data[44]
port 240 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 core_master_r_data[45]
port 241 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 core_master_r_data[46]
port 242 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 core_master_r_data[47]
port 243 nsew signal input
rlabel metal3 s 0 225768 800 225888 6 core_master_r_data[48]
port 244 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 core_master_r_data[49]
port 245 nsew signal input
rlabel metal3 s 279200 89088 280000 89208 6 core_master_r_data[4]
port 246 nsew signal input
rlabel metal2 s 229926 359200 229982 360000 6 core_master_r_data[50]
port 247 nsew signal input
rlabel metal2 s 119802 359200 119858 360000 6 core_master_r_data[51]
port 248 nsew signal input
rlabel metal3 s 279200 193808 280000 193928 6 core_master_r_data[52]
port 249 nsew signal input
rlabel metal2 s 153290 359200 153346 360000 6 core_master_r_data[53]
port 250 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 core_master_r_data[54]
port 251 nsew signal input
rlabel metal2 s 4526 359200 4582 360000 6 core_master_r_data[55]
port 252 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 core_master_r_data[56]
port 253 nsew signal input
rlabel metal3 s 279200 12248 280000 12368 6 core_master_r_data[57]
port 254 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 core_master_r_data[58]
port 255 nsew signal input
rlabel metal2 s 112718 359200 112774 360000 6 core_master_r_data[59]
port 256 nsew signal input
rlabel metal3 s 279200 42848 280000 42968 6 core_master_r_data[5]
port 257 nsew signal input
rlabel metal3 s 279200 335928 280000 336048 6 core_master_r_data[60]
port 258 nsew signal input
rlabel metal3 s 279200 20408 280000 20528 6 core_master_r_data[61]
port 259 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 core_master_r_data[62]
port 260 nsew signal input
rlabel metal2 s 219622 359200 219678 360000 6 core_master_r_data[63]
port 261 nsew signal input
rlabel metal2 s 153934 359200 153990 360000 6 core_master_r_data[6]
port 262 nsew signal input
rlabel metal2 s 150714 359200 150770 360000 6 core_master_r_data[7]
port 263 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 core_master_r_data[8]
port 264 nsew signal input
rlabel metal3 s 279200 140088 280000 140208 6 core_master_r_data[9]
port 265 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 core_master_r_id[0]
port 266 nsew signal input
rlabel metal2 s 9678 359200 9734 360000 6 core_master_r_id[1]
port 267 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 core_master_r_id[2]
port 268 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 core_master_r_id[3]
port 269 nsew signal input
rlabel metal3 s 0 346128 800 346248 6 core_master_r_id[4]
port 270 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 core_master_r_id[5]
port 271 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 core_master_r_id[6]
port 272 nsew signal input
rlabel metal3 s 0 239368 800 239488 6 core_master_r_id[7]
port 273 nsew signal input
rlabel metal2 s 242162 0 242218 800 6 core_master_r_id[8]
port 274 nsew signal input
rlabel metal3 s 279200 85008 280000 85128 6 core_master_r_id[9]
port 275 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 core_master_r_last
port 276 nsew signal input
rlabel metal3 s 279200 93168 280000 93288 6 core_master_r_ready
port 277 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 core_master_r_resp[0]
port 278 nsew signal input
rlabel metal3 s 279200 10888 280000 11008 6 core_master_r_resp[1]
port 279 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 core_master_r_user[-1]
port 280 nsew signal input
rlabel metal3 s 279200 144168 280000 144288 6 core_master_r_user[0]
port 281 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 core_master_r_valid
port 282 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 core_master_w_data[0]
port 283 nsew signal output
rlabel metal2 s 132038 359200 132094 360000 6 core_master_w_data[10]
port 284 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 core_master_w_data[11]
port 285 nsew signal output
rlabel metal3 s 0 176128 800 176248 6 core_master_w_data[12]
port 286 nsew signal output
rlabel metal3 s 279200 358368 280000 358488 6 core_master_w_data[13]
port 287 nsew signal output
rlabel metal3 s 0 318248 800 318368 6 core_master_w_data[14]
port 288 nsew signal output
rlabel metal2 s 198370 359200 198426 360000 6 core_master_w_data[15]
port 289 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 core_master_w_data[16]
port 290 nsew signal output
rlabel metal2 s 129462 359200 129518 360000 6 core_master_w_data[17]
port 291 nsew signal output
rlabel metal2 s 202234 0 202290 800 6 core_master_w_data[18]
port 292 nsew signal output
rlabel metal2 s 99838 359200 99894 360000 6 core_master_w_data[19]
port 293 nsew signal output
rlabel metal2 s 180338 359200 180394 360000 6 core_master_w_data[1]
port 294 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 core_master_w_data[20]
port 295 nsew signal output
rlabel metal3 s 279200 110168 280000 110288 6 core_master_w_data[21]
port 296 nsew signal output
rlabel metal3 s 0 285608 800 285728 6 core_master_w_data[22]
port 297 nsew signal output
rlabel metal3 s 279200 338648 280000 338768 6 core_master_w_data[23]
port 298 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 core_master_w_data[24]
port 299 nsew signal output
rlabel metal2 s 250534 359200 250590 360000 6 core_master_w_data[25]
port 300 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 core_master_w_data[26]
port 301 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 core_master_w_data[27]
port 302 nsew signal output
rlabel metal2 s 187422 359200 187478 360000 6 core_master_w_data[28]
port 303 nsew signal output
rlabel metal2 s 215758 359200 215814 360000 6 core_master_w_data[29]
port 304 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 core_master_w_data[2]
port 305 nsew signal output
rlabel metal3 s 279200 224408 280000 224528 6 core_master_w_data[30]
port 306 nsew signal output
rlabel metal3 s 0 191088 800 191208 6 core_master_w_data[31]
port 307 nsew signal output
rlabel metal3 s 0 181568 800 181688 6 core_master_w_data[32]
port 308 nsew signal output
rlabel metal3 s 279200 124448 280000 124568 6 core_master_w_data[33]
port 309 nsew signal output
rlabel metal3 s 279200 80928 280000 81048 6 core_master_w_data[34]
port 310 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 core_master_w_data[35]
port 311 nsew signal output
rlabel metal3 s 279200 64608 280000 64728 6 core_master_w_data[36]
port 312 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 core_master_w_data[37]
port 313 nsew signal output
rlabel metal2 s 65062 359200 65118 360000 6 core_master_w_data[38]
port 314 nsew signal output
rlabel metal2 s 114650 359200 114706 360000 6 core_master_w_data[39]
port 315 nsew signal output
rlabel metal3 s 279200 333888 280000 334008 6 core_master_w_data[3]
port 316 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 core_master_w_data[40]
port 317 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 core_master_w_data[41]
port 318 nsew signal output
rlabel metal3 s 0 315528 800 315648 6 core_master_w_data[42]
port 319 nsew signal output
rlabel metal3 s 279200 272688 280000 272808 6 core_master_w_data[43]
port 320 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 core_master_w_data[44]
port 321 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 core_master_w_data[45]
port 322 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 core_master_w_data[46]
port 323 nsew signal output
rlabel metal3 s 279200 99288 280000 99408 6 core_master_w_data[47]
port 324 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 core_master_w_data[48]
port 325 nsew signal output
rlabel metal3 s 0 241408 800 241528 6 core_master_w_data[49]
port 326 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 core_master_w_data[4]
port 327 nsew signal output
rlabel metal3 s 279200 18368 280000 18488 6 core_master_w_data[50]
port 328 nsew signal output
rlabel metal3 s 0 163888 800 164008 6 core_master_w_data[51]
port 329 nsew signal output
rlabel metal3 s 0 198568 800 198688 6 core_master_w_data[52]
port 330 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 core_master_w_data[53]
port 331 nsew signal output
rlabel metal2 s 184202 359200 184258 360000 6 core_master_w_data[54]
port 332 nsew signal output
rlabel metal3 s 0 339328 800 339448 6 core_master_w_data[55]
port 333 nsew signal output
rlabel metal2 s 63774 359200 63830 360000 6 core_master_w_data[56]
port 334 nsew signal output
rlabel metal3 s 279200 104048 280000 104168 6 core_master_w_data[57]
port 335 nsew signal output
rlabel metal3 s 279200 32648 280000 32768 6 core_master_w_data[58]
port 336 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 core_master_w_data[59]
port 337 nsew signal output
rlabel metal2 s 156510 359200 156566 360000 6 core_master_w_data[5]
port 338 nsew signal output
rlabel metal3 s 0 258408 800 258528 6 core_master_w_data[60]
port 339 nsew signal output
rlabel metal3 s 0 277448 800 277568 6 core_master_w_data[61]
port 340 nsew signal output
rlabel metal2 s 180338 0 180394 800 6 core_master_w_data[62]
port 341 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 core_master_w_data[63]
port 342 nsew signal output
rlabel metal3 s 279200 348168 280000 348288 6 core_master_w_data[6]
port 343 nsew signal output
rlabel metal2 s 255042 359200 255098 360000 6 core_master_w_data[7]
port 344 nsew signal output
rlabel metal3 s 279200 21768 280000 21888 6 core_master_w_data[8]
port 345 nsew signal output
rlabel metal3 s 0 170008 800 170128 6 core_master_w_data[9]
port 346 nsew signal output
rlabel metal2 s 208674 359200 208730 360000 6 core_master_w_last
port 347 nsew signal output
rlabel metal3 s 279200 91808 280000 91928 6 core_master_w_ready
port 348 nsew signal input
rlabel metal2 s 165526 359200 165582 360000 6 core_master_w_strb[0]
port 349 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 core_master_w_strb[1]
port 350 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 core_master_w_strb[2]
port 351 nsew signal output
rlabel metal3 s 279200 172728 280000 172848 6 core_master_w_strb[3]
port 352 nsew signal output
rlabel metal3 s 279200 176808 280000 176928 6 core_master_w_strb[4]
port 353 nsew signal output
rlabel metal3 s 279200 359048 280000 359168 6 core_master_w_strb[5]
port 354 nsew signal output
rlabel metal3 s 279200 125128 280000 125248 6 core_master_w_strb[6]
port 355 nsew signal output
rlabel metal3 s 279200 339328 280000 339448 6 core_master_w_strb[7]
port 356 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 core_master_w_user[-1]
port 357 nsew signal output
rlabel metal3 s 279200 55088 280000 55208 6 core_master_w_user[0]
port 358 nsew signal output
rlabel metal3 s 279200 169328 280000 169448 6 core_master_w_valid
port 359 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 data_slave_ar_addr[0]
port 360 nsew signal input
rlabel metal3 s 279200 223048 280000 223168 6 data_slave_ar_addr[10]
port 361 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 data_slave_ar_addr[11]
port 362 nsew signal input
rlabel metal2 s 271142 359200 271198 360000 6 data_slave_ar_addr[12]
port 363 nsew signal input
rlabel metal3 s 279200 39448 280000 39568 6 data_slave_ar_addr[13]
port 364 nsew signal input
rlabel metal3 s 279200 208768 280000 208888 6 data_slave_ar_addr[14]
port 365 nsew signal input
rlabel metal3 s 279200 181568 280000 181688 6 data_slave_ar_addr[15]
port 366 nsew signal input
rlabel metal3 s 0 227808 800 227928 6 data_slave_ar_addr[16]
port 367 nsew signal input
rlabel metal3 s 279200 309408 280000 309528 6 data_slave_ar_addr[17]
port 368 nsew signal input
rlabel metal3 s 279200 351568 280000 351688 6 data_slave_ar_addr[18]
port 369 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 data_slave_ar_addr[19]
port 370 nsew signal input
rlabel metal3 s 0 224408 800 224528 6 data_slave_ar_addr[1]
port 371 nsew signal input
rlabel metal2 s 97906 359200 97962 360000 6 data_slave_ar_addr[20]
port 372 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 data_slave_ar_addr[21]
port 373 nsew signal input
rlabel metal3 s 0 274728 800 274848 6 data_slave_ar_addr[22]
port 374 nsew signal input
rlabel metal2 s 268566 0 268622 800 6 data_slave_ar_addr[23]
port 375 nsew signal input
rlabel metal2 s 128174 359200 128230 360000 6 data_slave_ar_addr[24]
port 376 nsew signal input
rlabel metal2 s 258262 359200 258318 360000 6 data_slave_ar_addr[25]
port 377 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 data_slave_ar_addr[26]
port 378 nsew signal input
rlabel metal2 s 54758 359200 54814 360000 6 data_slave_ar_addr[27]
port 379 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 data_slave_ar_addr[28]
port 380 nsew signal input
rlabel metal3 s 279200 359728 280000 359848 6 data_slave_ar_addr[29]
port 381 nsew signal input
rlabel metal2 s 149426 359200 149482 360000 6 data_slave_ar_addr[2]
port 382 nsew signal input
rlabel metal3 s 0 232568 800 232688 6 data_slave_ar_addr[30]
port 383 nsew signal input
rlabel metal3 s 0 345448 800 345568 6 data_slave_ar_addr[31]
port 384 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 data_slave_ar_addr[3]
port 385 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 data_slave_ar_addr[4]
port 386 nsew signal input
rlabel metal3 s 279200 24488 280000 24608 6 data_slave_ar_addr[5]
port 387 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 data_slave_ar_addr[6]
port 388 nsew signal input
rlabel metal2 s 113362 359200 113418 360000 6 data_slave_ar_addr[7]
port 389 nsew signal input
rlabel metal2 s 142986 359200 143042 360000 6 data_slave_ar_addr[8]
port 390 nsew signal input
rlabel metal2 s 238298 359200 238354 360000 6 data_slave_ar_addr[9]
port 391 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 data_slave_ar_burst[0]
port 392 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 data_slave_ar_burst[1]
port 393 nsew signal input
rlabel metal3 s 279200 317568 280000 317688 6 data_slave_ar_cache[0]
port 394 nsew signal input
rlabel metal3 s 279200 11568 280000 11688 6 data_slave_ar_cache[1]
port 395 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 data_slave_ar_cache[2]
port 396 nsew signal input
rlabel metal2 s 168102 359200 168158 360000 6 data_slave_ar_cache[3]
port 397 nsew signal input
rlabel metal3 s 279200 82968 280000 83088 6 data_slave_ar_id[0]
port 398 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 data_slave_ar_id[1]
port 399 nsew signal input
rlabel metal3 s 279200 316208 280000 316328 6 data_slave_ar_id[2]
port 400 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 data_slave_ar_id[3]
port 401 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 data_slave_ar_id[4]
port 402 nsew signal input
rlabel metal3 s 279200 200608 280000 200728 6 data_slave_ar_id[5]
port 403 nsew signal input
rlabel metal3 s 279200 331848 280000 331968 6 data_slave_ar_id[6]
port 404 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 data_slave_ar_id[7]
port 405 nsew signal input
rlabel metal3 s 279200 37408 280000 37528 6 data_slave_ar_id[8]
port 406 nsew signal input
rlabel metal2 s 191930 359200 191986 360000 6 data_slave_ar_id[9]
port 407 nsew signal input
rlabel metal2 s 205454 359200 205510 360000 6 data_slave_ar_len[0]
port 408 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 data_slave_ar_len[1]
port 409 nsew signal input
rlabel metal2 s 132682 359200 132738 360000 6 data_slave_ar_len[2]
port 410 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 data_slave_ar_len[3]
port 411 nsew signal input
rlabel metal3 s 279200 346808 280000 346928 6 data_slave_ar_len[4]
port 412 nsew signal input
rlabel metal3 s 279200 265888 280000 266008 6 data_slave_ar_len[5]
port 413 nsew signal input
rlabel metal2 s 32218 359200 32274 360000 6 data_slave_ar_len[6]
port 414 nsew signal input
rlabel metal3 s 0 174768 800 174888 6 data_slave_ar_len[7]
port 415 nsew signal input
rlabel metal3 s 279200 152328 280000 152448 6 data_slave_ar_lock
port 416 nsew signal input
rlabel metal3 s 279200 36728 280000 36848 6 data_slave_ar_prot[0]
port 417 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 data_slave_ar_prot[1]
port 418 nsew signal input
rlabel metal3 s 0 356328 800 356448 6 data_slave_ar_prot[2]
port 419 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 data_slave_ar_qos[0]
port 420 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 data_slave_ar_qos[1]
port 421 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 data_slave_ar_qos[2]
port 422 nsew signal input
rlabel metal3 s 279200 330488 280000 330608 6 data_slave_ar_qos[3]
port 423 nsew signal input
rlabel metal3 s 0 351568 800 351688 6 data_slave_ar_ready
port 424 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 data_slave_ar_region[0]
port 425 nsew signal input
rlabel metal3 s 279200 133968 280000 134088 6 data_slave_ar_region[1]
port 426 nsew signal input
rlabel metal3 s 279200 49648 280000 49768 6 data_slave_ar_region[2]
port 427 nsew signal input
rlabel metal3 s 0 307368 800 307488 6 data_slave_ar_region[3]
port 428 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 data_slave_ar_size[0]
port 429 nsew signal input
rlabel metal3 s 279200 270648 280000 270768 6 data_slave_ar_size[1]
port 430 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 data_slave_ar_size[2]
port 431 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 data_slave_ar_user[-1]
port 432 nsew signal input
rlabel metal3 s 0 187008 800 187128 6 data_slave_ar_user[0]
port 433 nsew signal input
rlabel metal2 s 184846 0 184902 800 6 data_slave_ar_valid
port 434 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 data_slave_aw_addr[0]
port 435 nsew signal input
rlabel metal3 s 279200 235288 280000 235408 6 data_slave_aw_addr[10]
port 436 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 data_slave_aw_addr[11]
port 437 nsew signal input
rlabel metal3 s 0 221008 800 221128 6 data_slave_aw_addr[12]
port 438 nsew signal input
rlabel metal2 s 224130 359200 224186 360000 6 data_slave_aw_addr[13]
port 439 nsew signal input
rlabel metal2 s 82450 359200 82506 360000 6 data_slave_aw_addr[14]
port 440 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 data_slave_aw_addr[15]
port 441 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 data_slave_aw_addr[16]
port 442 nsew signal input
rlabel metal3 s 0 296488 800 296608 6 data_slave_aw_addr[17]
port 443 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 data_slave_aw_addr[18]
port 444 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 data_slave_aw_addr[19]
port 445 nsew signal input
rlabel metal2 s 175186 359200 175242 360000 6 data_slave_aw_addr[1]
port 446 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 data_slave_aw_addr[20]
port 447 nsew signal input
rlabel metal3 s 0 148928 800 149048 6 data_slave_aw_addr[21]
port 448 nsew signal input
rlabel metal3 s 279200 228488 280000 228608 6 data_slave_aw_addr[22]
port 449 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 data_slave_aw_addr[23]
port 450 nsew signal input
rlabel metal3 s 0 226448 800 226568 6 data_slave_aw_addr[24]
port 451 nsew signal input
rlabel metal2 s 66994 359200 67050 360000 6 data_slave_aw_addr[25]
port 452 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 data_slave_aw_addr[26]
port 453 nsew signal input
rlabel metal3 s 0 195848 800 195968 6 data_slave_aw_addr[27]
port 454 nsew signal input
rlabel metal3 s 0 338648 800 338768 6 data_slave_aw_addr[28]
port 455 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 data_slave_aw_addr[29]
port 456 nsew signal input
rlabel metal3 s 279200 4768 280000 4888 6 data_slave_aw_addr[2]
port 457 nsew signal input
rlabel metal2 s 155222 359200 155278 360000 6 data_slave_aw_addr[30]
port 458 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 data_slave_aw_addr[31]
port 459 nsew signal input
rlabel metal2 s 86958 359200 87014 360000 6 data_slave_aw_addr[3]
port 460 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 data_slave_aw_addr[4]
port 461 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 data_slave_aw_addr[5]
port 462 nsew signal input
rlabel metal2 s 273074 359200 273130 360000 6 data_slave_aw_addr[6]
port 463 nsew signal input
rlabel metal3 s 279200 19728 280000 19848 6 data_slave_aw_addr[7]
port 464 nsew signal input
rlabel metal3 s 279200 138048 280000 138168 6 data_slave_aw_addr[8]
port 465 nsew signal input
rlabel metal2 s 238942 0 238998 800 6 data_slave_aw_addr[9]
port 466 nsew signal input
rlabel metal3 s 0 243448 800 243568 6 data_slave_aw_burst[0]
port 467 nsew signal input
rlabel metal3 s 0 144848 800 144968 6 data_slave_aw_burst[1]
port 468 nsew signal input
rlabel metal3 s 279200 332528 280000 332648 6 data_slave_aw_cache[0]
port 469 nsew signal input
rlabel metal3 s 0 175448 800 175568 6 data_slave_aw_cache[1]
port 470 nsew signal input
rlabel metal3 s 279200 187688 280000 187808 6 data_slave_aw_cache[2]
port 471 nsew signal input
rlabel metal3 s 0 359048 800 359168 6 data_slave_aw_cache[3]
port 472 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 data_slave_aw_id[0]
port 473 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 data_slave_aw_id[1]
port 474 nsew signal input
rlabel metal3 s 279200 297168 280000 297288 6 data_slave_aw_id[2]
port 475 nsew signal input
rlabel metal3 s 0 201288 800 201408 6 data_slave_aw_id[3]
port 476 nsew signal input
rlabel metal3 s 0 304648 800 304768 6 data_slave_aw_id[4]
port 477 nsew signal input
rlabel metal3 s 279200 242088 280000 242208 6 data_slave_aw_id[5]
port 478 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 data_slave_aw_id[6]
port 479 nsew signal input
rlabel metal2 s 83738 359200 83794 360000 6 data_slave_aw_id[7]
port 480 nsew signal input
rlabel metal3 s 279200 41488 280000 41608 6 data_slave_aw_id[8]
port 481 nsew signal input
rlabel metal2 s 71502 359200 71558 360000 6 data_slave_aw_id[9]
port 482 nsew signal input
rlabel metal3 s 279200 133288 280000 133408 6 data_slave_aw_len[0]
port 483 nsew signal input
rlabel metal3 s 279200 106088 280000 106208 6 data_slave_aw_len[1]
port 484 nsew signal input
rlabel metal3 s 0 331848 800 331968 6 data_slave_aw_len[2]
port 485 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 data_slave_aw_len[3]
port 486 nsew signal input
rlabel metal3 s 279200 278808 280000 278928 6 data_slave_aw_len[4]
port 487 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 data_slave_aw_len[5]
port 488 nsew signal input
rlabel metal2 s 69570 359200 69626 360000 6 data_slave_aw_len[6]
port 489 nsew signal input
rlabel metal3 s 0 335928 800 336048 6 data_slave_aw_len[7]
port 490 nsew signal input
rlabel metal2 s 1306 359200 1362 360000 6 data_slave_aw_lock
port 491 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 data_slave_aw_prot[0]
port 492 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 data_slave_aw_prot[1]
port 493 nsew signal input
rlabel metal2 s 662 359200 718 360000 6 data_slave_aw_prot[2]
port 494 nsew signal input
rlabel metal3 s 279200 92488 280000 92608 6 data_slave_aw_qos[0]
port 495 nsew signal input
rlabel metal3 s 279200 50328 280000 50448 6 data_slave_aw_qos[1]
port 496 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 data_slave_aw_qos[2]
port 497 nsew signal input
rlabel metal3 s 279200 298528 280000 298648 6 data_slave_aw_qos[3]
port 498 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 data_slave_aw_ready
port 499 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 data_slave_aw_region[0]
port 500 nsew signal input
rlabel metal3 s 279200 303288 280000 303408 6 data_slave_aw_region[1]
port 501 nsew signal input
rlabel metal3 s 279200 343408 280000 343528 6 data_slave_aw_region[2]
port 502 nsew signal input
rlabel metal3 s 0 169328 800 169448 6 data_slave_aw_region[3]
port 503 nsew signal input
rlabel metal3 s 0 215568 800 215688 6 data_slave_aw_size[0]
port 504 nsew signal input
rlabel metal3 s 0 193128 800 193248 6 data_slave_aw_size[1]
port 505 nsew signal input
rlabel metal3 s 0 306688 800 306808 6 data_slave_aw_size[2]
port 506 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 data_slave_aw_user[-1]
port 507 nsew signal input
rlabel metal2 s 223486 359200 223542 360000 6 data_slave_aw_user[0]
port 508 nsew signal input
rlabel metal3 s 279200 261808 280000 261928 6 data_slave_aw_valid
port 509 nsew signal input
rlabel metal3 s 279200 167968 280000 168088 6 data_slave_b_id[0]
port 510 nsew signal output
rlabel metal3 s 279200 306008 280000 306128 6 data_slave_b_id[1]
port 511 nsew signal output
rlabel metal2 s 29642 359200 29698 360000 6 data_slave_b_id[2]
port 512 nsew signal output
rlabel metal3 s 0 344088 800 344208 6 data_slave_b_id[3]
port 513 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 data_slave_b_id[4]
port 514 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 data_slave_b_id[5]
port 515 nsew signal output
rlabel metal3 s 0 282208 800 282328 6 data_slave_b_id[6]
port 516 nsew signal output
rlabel metal3 s 279200 130568 280000 130688 6 data_slave_b_id[7]
port 517 nsew signal output
rlabel metal3 s 279200 352248 280000 352368 6 data_slave_b_id[8]
port 518 nsew signal output
rlabel metal3 s 0 276768 800 276888 6 data_slave_b_id[9]
port 519 nsew signal output
rlabel metal2 s 143630 359200 143686 360000 6 data_slave_b_ready
port 520 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 data_slave_b_resp[0]
port 521 nsew signal output
rlabel metal2 s 195150 359200 195206 360000 6 data_slave_b_resp[1]
port 522 nsew signal output
rlabel metal3 s 279200 102008 280000 102128 6 data_slave_b_user[-1]
port 523 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 data_slave_b_user[0]
port 524 nsew signal output
rlabel metal3 s 0 183608 800 183728 6 data_slave_b_valid
port 525 nsew signal output
rlabel metal2 s 110786 359200 110842 360000 6 data_slave_r_data[0]
port 526 nsew signal output
rlabel metal3 s 279200 240048 280000 240168 6 data_slave_r_data[10]
port 527 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 data_slave_r_data[11]
port 528 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 data_slave_r_data[12]
port 529 nsew signal output
rlabel metal2 s 276938 359200 276994 360000 6 data_slave_r_data[13]
port 530 nsew signal output
rlabel metal3 s 0 279488 800 279608 6 data_slave_r_data[14]
port 531 nsew signal output
rlabel metal2 s 242806 359200 242862 360000 6 data_slave_r_data[15]
port 532 nsew signal output
rlabel metal3 s 279200 97928 280000 98048 6 data_slave_r_data[16]
port 533 nsew signal output
rlabel metal3 s 0 214208 800 214328 6 data_slave_r_data[17]
port 534 nsew signal output
rlabel metal2 s 197726 0 197782 800 6 data_slave_r_data[18]
port 535 nsew signal output
rlabel metal2 s 182914 0 182970 800 6 data_slave_r_data[19]
port 536 nsew signal output
rlabel metal3 s 0 344768 800 344888 6 data_slave_r_data[1]
port 537 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 data_slave_r_data[20]
port 538 nsew signal output
rlabel metal2 s 3238 359200 3294 360000 6 data_slave_r_data[21]
port 539 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 data_slave_r_data[22]
port 540 nsew signal output
rlabel metal2 s 270498 0 270554 800 6 data_slave_r_data[23]
port 541 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 data_slave_r_data[24]
port 542 nsew signal output
rlabel metal2 s 110142 359200 110198 360000 6 data_slave_r_data[25]
port 543 nsew signal output
rlabel metal2 s 59266 359200 59322 360000 6 data_slave_r_data[26]
port 544 nsew signal output
rlabel metal3 s 0 262488 800 262608 6 data_slave_r_data[27]
port 545 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 data_slave_r_data[28]
port 546 nsew signal output
rlabel metal2 s 92110 359200 92166 360000 6 data_slave_r_data[29]
port 547 nsew signal output
rlabel metal3 s 279200 195848 280000 195968 6 data_slave_r_data[2]
port 548 nsew signal output
rlabel metal3 s 279200 149608 280000 149728 6 data_slave_r_data[30]
port 549 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 data_slave_r_data[31]
port 550 nsew signal output
rlabel metal2 s 181626 0 181682 800 6 data_slave_r_data[32]
port 551 nsew signal output
rlabel metal3 s 0 320288 800 320408 6 data_slave_r_data[33]
port 552 nsew signal output
rlabel metal2 s 213826 0 213882 800 6 data_slave_r_data[34]
port 553 nsew signal output
rlabel metal3 s 279200 217608 280000 217728 6 data_slave_r_data[35]
port 554 nsew signal output
rlabel metal3 s 0 352928 800 353048 6 data_slave_r_data[36]
port 555 nsew signal output
rlabel metal3 s 279200 191768 280000 191888 6 data_slave_r_data[37]
port 556 nsew signal output
rlabel metal2 s 231858 0 231914 800 6 data_slave_r_data[38]
port 557 nsew signal output
rlabel metal2 s 253754 0 253810 800 6 data_slave_r_data[39]
port 558 nsew signal output
rlabel metal3 s 0 286288 800 286408 6 data_slave_r_data[3]
port 559 nsew signal output
rlabel metal2 s 144918 359200 144974 360000 6 data_slave_r_data[40]
port 560 nsew signal output
rlabel metal2 s 18 359200 74 360000 6 data_slave_r_data[41]
port 561 nsew signal output
rlabel metal2 s 107566 359200 107622 360000 6 data_slave_r_data[42]
port 562 nsew signal output
rlabel metal2 s 214470 359200 214526 360000 6 data_slave_r_data[43]
port 563 nsew signal output
rlabel metal3 s 279200 123768 280000 123888 6 data_slave_r_data[44]
port 564 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 data_slave_r_data[45]
port 565 nsew signal output
rlabel metal3 s 0 213528 800 213648 6 data_slave_r_data[46]
port 566 nsew signal output
rlabel metal2 s 196438 359200 196494 360000 6 data_slave_r_data[47]
port 567 nsew signal output
rlabel metal3 s 279200 331168 280000 331288 6 data_slave_r_data[48]
port 568 nsew signal output
rlabel metal3 s 279200 36048 280000 36168 6 data_slave_r_data[49]
port 569 nsew signal output
rlabel metal2 s 201590 0 201646 800 6 data_slave_r_data[4]
port 570 nsew signal output
rlabel metal3 s 0 264528 800 264648 6 data_slave_r_data[50]
port 571 nsew signal output
rlabel metal3 s 279200 146208 280000 146328 6 data_slave_r_data[51]
port 572 nsew signal output
rlabel metal3 s 0 322328 800 322448 6 data_slave_r_data[52]
port 573 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 data_slave_r_data[53]
port 574 nsew signal output
rlabel metal3 s 279200 146888 280000 147008 6 data_slave_r_data[54]
port 575 nsew signal output
rlabel metal3 s 279200 119008 280000 119128 6 data_slave_r_data[55]
port 576 nsew signal output
rlabel metal3 s 0 237328 800 237448 6 data_slave_r_data[56]
port 577 nsew signal output
rlabel metal3 s 279200 82288 280000 82408 6 data_slave_r_data[57]
port 578 nsew signal output
rlabel metal2 s 50250 359200 50306 360000 6 data_slave_r_data[58]
port 579 nsew signal output
rlabel metal2 s 19338 359200 19394 360000 6 data_slave_r_data[59]
port 580 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 data_slave_r_data[5]
port 581 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 data_slave_r_data[60]
port 582 nsew signal output
rlabel metal3 s 0 269288 800 269408 6 data_slave_r_data[61]
port 583 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 data_slave_r_data[62]
port 584 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 data_slave_r_data[63]
port 585 nsew signal output
rlabel metal2 s 216402 0 216458 800 6 data_slave_r_data[6]
port 586 nsew signal output
rlabel metal2 s 248602 359200 248658 360000 6 data_slave_r_data[7]
port 587 nsew signal output
rlabel metal2 s 267278 359200 267334 360000 6 data_slave_r_data[8]
port 588 nsew signal output
rlabel metal3 s 279200 290368 280000 290488 6 data_slave_r_data[9]
port 589 nsew signal output
rlabel metal3 s 279200 108808 280000 108928 6 data_slave_r_id[0]
port 590 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 data_slave_r_id[1]
port 591 nsew signal output
rlabel metal3 s 279200 225768 280000 225888 6 data_slave_r_id[2]
port 592 nsew signal output
rlabel metal3 s 279200 255688 280000 255808 6 data_slave_r_id[3]
port 593 nsew signal output
rlabel metal2 s 166814 0 166870 800 6 data_slave_r_id[4]
port 594 nsew signal output
rlabel metal2 s 271786 0 271842 800 6 data_slave_r_id[5]
port 595 nsew signal output
rlabel metal2 s 6458 359200 6514 360000 6 data_slave_r_id[6]
port 596 nsew signal output
rlabel metal3 s 0 214888 800 215008 6 data_slave_r_id[7]
port 597 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 data_slave_r_id[8]
port 598 nsew signal output
rlabel metal3 s 279200 333208 280000 333328 6 data_slave_r_id[9]
port 599 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 data_slave_r_last
port 600 nsew signal output
rlabel metal2 s 265990 0 266046 800 6 data_slave_r_ready
port 601 nsew signal input
rlabel metal2 s 276294 359200 276350 360000 6 data_slave_r_resp[0]
port 602 nsew signal output
rlabel metal3 s 279200 117648 280000 117768 6 data_slave_r_resp[1]
port 603 nsew signal output
rlabel metal2 s 179694 359200 179750 360000 6 data_slave_r_user[-1]
port 604 nsew signal output
rlabel metal3 s 279200 74128 280000 74248 6 data_slave_r_user[0]
port 605 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 data_slave_r_valid
port 606 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 data_slave_w_data[0]
port 607 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 data_slave_w_data[10]
port 608 nsew signal input
rlabel metal2 s 157154 359200 157210 360000 6 data_slave_w_data[11]
port 609 nsew signal input
rlabel metal2 s 246670 359200 246726 360000 6 data_slave_w_data[12]
port 610 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 data_slave_w_data[13]
port 611 nsew signal input
rlabel metal3 s 0 261128 800 261248 6 data_slave_w_data[14]
port 612 nsew signal input
rlabel metal2 s 88246 359200 88302 360000 6 data_slave_w_data[15]
port 613 nsew signal input
rlabel metal3 s 0 281528 800 281648 6 data_slave_w_data[16]
port 614 nsew signal input
rlabel metal2 s 137834 359200 137890 360000 6 data_slave_w_data[17]
port 615 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 data_slave_w_data[18]
port 616 nsew signal input
rlabel metal3 s 279200 74808 280000 74928 6 data_slave_w_data[19]
port 617 nsew signal input
rlabel metal3 s 279200 272008 280000 272128 6 data_slave_w_data[1]
port 618 nsew signal input
rlabel metal3 s 0 291728 800 291848 6 data_slave_w_data[20]
port 619 nsew signal input
rlabel metal2 s 7102 359200 7158 360000 6 data_slave_w_data[21]
port 620 nsew signal input
rlabel metal3 s 279200 161168 280000 161288 6 data_slave_w_data[22]
port 621 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 data_slave_w_data[23]
port 622 nsew signal input
rlabel metal2 s 67638 359200 67694 360000 6 data_slave_w_data[24]
port 623 nsew signal input
rlabel metal3 s 279200 284248 280000 284368 6 data_slave_w_data[25]
port 624 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 data_slave_w_data[26]
port 625 nsew signal input
rlabel metal3 s 0 199928 800 200048 6 data_slave_w_data[27]
port 626 nsew signal input
rlabel metal3 s 279200 314168 280000 314288 6 data_slave_w_data[28]
port 627 nsew signal input
rlabel metal2 s 105634 359200 105690 360000 6 data_slave_w_data[29]
port 628 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 data_slave_w_data[2]
port 629 nsew signal input
rlabel metal2 s 22558 359200 22614 360000 6 data_slave_w_data[30]
port 630 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 data_slave_w_data[31]
port 631 nsew signal input
rlabel metal3 s 279200 26528 280000 26648 6 data_slave_w_data[32]
port 632 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 data_slave_w_data[33]
port 633 nsew signal input
rlabel metal3 s 0 335248 800 335368 6 data_slave_w_data[34]
port 634 nsew signal input
rlabel metal3 s 0 138048 800 138168 6 data_slave_w_data[35]
port 635 nsew signal input
rlabel metal2 s 57334 359200 57390 360000 6 data_slave_w_data[36]
port 636 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 data_slave_w_data[37]
port 637 nsew signal input
rlabel metal3 s 279200 3408 280000 3528 6 data_slave_w_data[38]
port 638 nsew signal input
rlabel metal2 s 21914 359200 21970 360000 6 data_slave_w_data[39]
port 639 nsew signal input
rlabel metal3 s 279200 29928 280000 30048 6 data_slave_w_data[3]
port 640 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 data_slave_w_data[40]
port 641 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 data_slave_w_data[41]
port 642 nsew signal input
rlabel metal2 s 211894 359200 211950 360000 6 data_slave_w_data[42]
port 643 nsew signal input
rlabel metal2 s 177762 359200 177818 360000 6 data_slave_w_data[43]
port 644 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 data_slave_w_data[44]
port 645 nsew signal input
rlabel metal3 s 279200 172048 280000 172168 6 data_slave_w_data[45]
port 646 nsew signal input
rlabel metal2 s 34794 359200 34850 360000 6 data_slave_w_data[46]
port 647 nsew signal input
rlabel metal2 s 58622 359200 58678 360000 6 data_slave_w_data[47]
port 648 nsew signal input
rlabel metal3 s 0 313488 800 313608 6 data_slave_w_data[48]
port 649 nsew signal input
rlabel metal2 s 209962 0 210018 800 6 data_slave_w_data[49]
port 650 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 data_slave_w_data[4]
port 651 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 data_slave_w_data[50]
port 652 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 data_slave_w_data[51]
port 653 nsew signal input
rlabel metal3 s 279200 125808 280000 125928 6 data_slave_w_data[52]
port 654 nsew signal input
rlabel metal3 s 279200 80248 280000 80368 6 data_slave_w_data[53]
port 655 nsew signal input
rlabel metal2 s 135902 359200 135958 360000 6 data_slave_w_data[54]
port 656 nsew signal input
rlabel metal3 s 279200 66648 280000 66768 6 data_slave_w_data[55]
port 657 nsew signal input
rlabel metal3 s 0 129888 800 130008 6 data_slave_w_data[56]
port 658 nsew signal input
rlabel metal2 s 265346 359200 265402 360000 6 data_slave_w_data[57]
port 659 nsew signal input
rlabel metal2 s 263414 0 263470 800 6 data_slave_w_data[58]
port 660 nsew signal input
rlabel metal2 s 133970 359200 134026 360000 6 data_slave_w_data[59]
port 661 nsew signal input
rlabel metal3 s 279200 204688 280000 204808 6 data_slave_w_data[5]
port 662 nsew signal input
rlabel metal2 s 146206 359200 146262 360000 6 data_slave_w_data[60]
port 663 nsew signal input
rlabel metal2 s 201590 359200 201646 360000 6 data_slave_w_data[61]
port 664 nsew signal input
rlabel metal2 s 244094 359200 244150 360000 6 data_slave_w_data[62]
port 665 nsew signal input
rlabel metal3 s 279200 114928 280000 115048 6 data_slave_w_data[63]
port 666 nsew signal input
rlabel metal2 s 116582 359200 116638 360000 6 data_slave_w_data[6]
port 667 nsew signal input
rlabel metal3 s 279200 142808 280000 142928 6 data_slave_w_data[7]
port 668 nsew signal input
rlabel metal2 s 164882 359200 164938 360000 6 data_slave_w_data[8]
port 669 nsew signal input
rlabel metal3 s 0 299888 800 300008 6 data_slave_w_data[9]
port 670 nsew signal input
rlabel metal3 s 279200 300568 280000 300688 6 data_slave_w_last
port 671 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 data_slave_w_ready
port 672 nsew signal output
rlabel metal3 s 279200 325048 280000 325168 6 data_slave_w_strb[0]
port 673 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 data_slave_w_strb[1]
port 674 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 data_slave_w_strb[2]
port 675 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 data_slave_w_strb[3]
port 676 nsew signal input
rlabel metal2 s 77942 359200 77998 360000 6 data_slave_w_strb[4]
port 677 nsew signal input
rlabel metal3 s 279200 136008 280000 136128 6 data_slave_w_strb[5]
port 678 nsew signal input
rlabel metal2 s 39946 359200 40002 360000 6 data_slave_w_strb[6]
port 679 nsew signal input
rlabel metal3 s 279200 138728 280000 138848 6 data_slave_w_strb[7]
port 680 nsew signal input
rlabel metal3 s 279200 132608 280000 132728 6 data_slave_w_user[-1]
port 681 nsew signal input
rlabel metal3 s 279200 206728 280000 206848 6 data_slave_w_user[0]
port 682 nsew signal input
rlabel metal2 s 159730 359200 159786 360000 6 data_slave_w_valid
port 683 nsew signal input
rlabel metal3 s 279200 262488 280000 262608 6 dbg_master_ar_addr[0]
port 684 nsew signal output
rlabel metal3 s 0 261808 800 261928 6 dbg_master_ar_addr[10]
port 685 nsew signal output
rlabel metal3 s 279200 13608 280000 13728 6 dbg_master_ar_addr[11]
port 686 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 dbg_master_ar_addr[12]
port 687 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 dbg_master_ar_addr[13]
port 688 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 dbg_master_ar_addr[14]
port 689 nsew signal output
rlabel metal3 s 279200 278128 280000 278248 6 dbg_master_ar_addr[15]
port 690 nsew signal output
rlabel metal2 s 238298 0 238354 800 6 dbg_master_ar_addr[16]
port 691 nsew signal output
rlabel metal3 s 279200 129888 280000 130008 6 dbg_master_ar_addr[17]
port 692 nsew signal output
rlabel metal3 s 279200 112888 280000 113008 6 dbg_master_ar_addr[18]
port 693 nsew signal output
rlabel metal2 s 187422 0 187478 800 6 dbg_master_ar_addr[19]
port 694 nsew signal output
rlabel metal2 s 204810 0 204866 800 6 dbg_master_ar_addr[1]
port 695 nsew signal output
rlabel metal2 s 146850 359200 146906 360000 6 dbg_master_ar_addr[20]
port 696 nsew signal output
rlabel metal2 s 206098 359200 206154 360000 6 dbg_master_ar_addr[21]
port 697 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 dbg_master_ar_addr[22]
port 698 nsew signal output
rlabel metal2 s 270498 359200 270554 360000 6 dbg_master_ar_addr[23]
port 699 nsew signal output
rlabel metal2 s 195794 359200 195850 360000 6 dbg_master_ar_addr[24]
port 700 nsew signal output
rlabel metal3 s 279200 170688 280000 170808 6 dbg_master_ar_addr[25]
port 701 nsew signal output
rlabel metal3 s 0 148248 800 148368 6 dbg_master_ar_addr[26]
port 702 nsew signal output
rlabel metal2 s 186134 359200 186190 360000 6 dbg_master_ar_addr[27]
port 703 nsew signal output
rlabel metal3 s 279200 288328 280000 288448 6 dbg_master_ar_addr[28]
port 704 nsew signal output
rlabel metal3 s 279200 196528 280000 196648 6 dbg_master_ar_addr[29]
port 705 nsew signal output
rlabel metal3 s 279200 293768 280000 293888 6 dbg_master_ar_addr[2]
port 706 nsew signal output
rlabel metal2 s 68926 359200 68982 360000 6 dbg_master_ar_addr[30]
port 707 nsew signal output
rlabel metal2 s 50894 359200 50950 360000 6 dbg_master_ar_addr[31]
port 708 nsew signal output
rlabel metal2 s 211894 0 211950 800 6 dbg_master_ar_addr[3]
port 709 nsew signal output
rlabel metal3 s 279200 216248 280000 216368 6 dbg_master_ar_addr[4]
port 710 nsew signal output
rlabel metal3 s 0 245488 800 245608 6 dbg_master_ar_addr[5]
port 711 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 dbg_master_ar_addr[6]
port 712 nsew signal output
rlabel metal2 s 2594 359200 2650 360000 6 dbg_master_ar_addr[7]
port 713 nsew signal output
rlabel metal3 s 279200 197888 280000 198008 6 dbg_master_ar_addr[8]
port 714 nsew signal output
rlabel metal2 s 235078 359200 235134 360000 6 dbg_master_ar_addr[9]
port 715 nsew signal output
rlabel metal3 s 0 165928 800 166048 6 dbg_master_ar_burst[0]
port 716 nsew signal output
rlabel metal3 s 279200 260448 280000 260568 6 dbg_master_ar_burst[1]
port 717 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 dbg_master_ar_cache[0]
port 718 nsew signal output
rlabel metal3 s 0 217608 800 217728 6 dbg_master_ar_cache[1]
port 719 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 dbg_master_ar_cache[2]
port 720 nsew signal output
rlabel metal2 s 212538 0 212594 800 6 dbg_master_ar_cache[3]
port 721 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 dbg_master_ar_id[0]
port 722 nsew signal output
rlabel metal2 s 108854 359200 108910 360000 6 dbg_master_ar_id[1]
port 723 nsew signal output
rlabel metal2 s 278870 0 278926 800 6 dbg_master_ar_id[2]
port 724 nsew signal output
rlabel metal3 s 0 326408 800 326528 6 dbg_master_ar_id[3]
port 725 nsew signal output
rlabel metal3 s 279200 88408 280000 88528 6 dbg_master_ar_id[4]
port 726 nsew signal output
rlabel metal2 s 227350 359200 227406 360000 6 dbg_master_ar_id[5]
port 727 nsew signal output
rlabel metal3 s 0 216248 800 216368 6 dbg_master_ar_id[6]
port 728 nsew signal output
rlabel metal3 s 279200 310768 280000 310888 6 dbg_master_ar_id[7]
port 729 nsew signal output
rlabel metal3 s 279200 244808 280000 244928 6 dbg_master_ar_id[8]
port 730 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 dbg_master_ar_id[9]
port 731 nsew signal output
rlabel metal3 s 0 255688 800 255808 6 dbg_master_ar_len[0]
port 732 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 dbg_master_ar_len[1]
port 733 nsew signal output
rlabel metal3 s 279200 29248 280000 29368 6 dbg_master_ar_len[2]
port 734 nsew signal output
rlabel metal2 s 216402 359200 216458 360000 6 dbg_master_ar_len[3]
port 735 nsew signal output
rlabel metal2 s 119158 359200 119214 360000 6 dbg_master_ar_len[4]
port 736 nsew signal output
rlabel metal2 s 77298 359200 77354 360000 6 dbg_master_ar_len[5]
port 737 nsew signal output
rlabel metal3 s 0 235968 800 236088 6 dbg_master_ar_len[6]
port 738 nsew signal output
rlabel metal3 s 0 155728 800 155848 6 dbg_master_ar_len[7]
port 739 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 dbg_master_ar_lock
port 740 nsew signal output
rlabel metal3 s 0 289688 800 289808 6 dbg_master_ar_prot[0]
port 741 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 dbg_master_ar_prot[1]
port 742 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 dbg_master_ar_prot[2]
port 743 nsew signal output
rlabel metal2 s 93398 359200 93454 360000 6 dbg_master_ar_qos[0]
port 744 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 dbg_master_ar_qos[1]
port 745 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 dbg_master_ar_qos[2]
port 746 nsew signal output
rlabel metal2 s 211250 0 211306 800 6 dbg_master_ar_qos[3]
port 747 nsew signal output
rlabel metal3 s 279200 209448 280000 209568 6 dbg_master_ar_ready
port 748 nsew signal input
rlabel metal2 s 141698 359200 141754 360000 6 dbg_master_ar_region[0]
port 749 nsew signal output
rlabel metal2 s 227994 359200 228050 360000 6 dbg_master_ar_region[1]
port 750 nsew signal output
rlabel metal3 s 0 223728 800 223848 6 dbg_master_ar_region[2]
port 751 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 dbg_master_ar_region[3]
port 752 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 dbg_master_ar_size[0]
port 753 nsew signal output
rlabel metal2 s 76654 359200 76710 360000 6 dbg_master_ar_size[1]
port 754 nsew signal output
rlabel metal2 s 126242 359200 126298 360000 6 dbg_master_ar_size[2]
port 755 nsew signal output
rlabel metal2 s 43810 359200 43866 360000 6 dbg_master_ar_user[-1]
port 756 nsew signal output
rlabel metal2 s 208674 0 208730 800 6 dbg_master_ar_user[0]
port 757 nsew signal output
rlabel metal2 s 103702 359200 103758 360000 6 dbg_master_ar_valid
port 758 nsew signal output
rlabel metal2 s 13542 359200 13598 360000 6 dbg_master_aw_addr[0]
port 759 nsew signal output
rlabel metal3 s 279200 65968 280000 66088 6 dbg_master_aw_addr[10]
port 760 nsew signal output
rlabel metal3 s 279200 337968 280000 338088 6 dbg_master_aw_addr[11]
port 761 nsew signal output
rlabel metal2 s 80518 359200 80574 360000 6 dbg_master_aw_addr[12]
port 762 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 dbg_master_aw_addr[13]
port 763 nsew signal output
rlabel metal3 s 279200 107448 280000 107568 6 dbg_master_aw_addr[14]
port 764 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 dbg_master_aw_addr[15]
port 765 nsew signal output
rlabel metal3 s 0 182248 800 182368 6 dbg_master_aw_addr[16]
port 766 nsew signal output
rlabel metal2 s 136546 359200 136602 360000 6 dbg_master_aw_addr[17]
port 767 nsew signal output
rlabel metal3 s 279200 323688 280000 323808 6 dbg_master_aw_addr[18]
port 768 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 dbg_master_aw_addr[19]
port 769 nsew signal output
rlabel metal3 s 279200 357688 280000 357808 6 dbg_master_aw_addr[1]
port 770 nsew signal output
rlabel metal3 s 279200 111528 280000 111648 6 dbg_master_aw_addr[20]
port 771 nsew signal output
rlabel metal2 s 45098 359200 45154 360000 6 dbg_master_aw_addr[21]
port 772 nsew signal output
rlabel metal2 s 140410 0 140466 800 6 dbg_master_aw_addr[22]
port 773 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 dbg_master_aw_addr[23]
port 774 nsew signal output
rlabel metal3 s 279200 245488 280000 245608 6 dbg_master_aw_addr[24]
port 775 nsew signal output
rlabel metal2 s 247314 359200 247370 360000 6 dbg_master_aw_addr[25]
port 776 nsew signal output
rlabel metal3 s 279200 249568 280000 249688 6 dbg_master_aw_addr[26]
port 777 nsew signal output
rlabel metal3 s 0 123088 800 123208 6 dbg_master_aw_addr[27]
port 778 nsew signal output
rlabel metal2 s 130750 359200 130806 360000 6 dbg_master_aw_addr[28]
port 779 nsew signal output
rlabel metal3 s 0 233248 800 233368 6 dbg_master_aw_addr[29]
port 780 nsew signal output
rlabel metal3 s 0 298528 800 298648 6 dbg_master_aw_addr[2]
port 781 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 dbg_master_aw_addr[30]
port 782 nsew signal output
rlabel metal2 s 268566 359200 268622 360000 6 dbg_master_aw_addr[31]
port 783 nsew signal output
rlabel metal2 s 239586 359200 239642 360000 6 dbg_master_aw_addr[3]
port 784 nsew signal output
rlabel metal3 s 279200 310088 280000 310208 6 dbg_master_aw_addr[4]
port 785 nsew signal output
rlabel metal3 s 0 340008 800 340128 6 dbg_master_aw_addr[5]
port 786 nsew signal output
rlabel metal3 s 279200 183608 280000 183728 6 dbg_master_aw_addr[6]
port 787 nsew signal output
rlabel metal3 s 279200 350208 280000 350328 6 dbg_master_aw_addr[7]
port 788 nsew signal output
rlabel metal2 s 247314 0 247370 800 6 dbg_master_aw_addr[8]
port 789 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 dbg_master_aw_addr[9]
port 790 nsew signal output
rlabel metal3 s 279200 21088 280000 21208 6 dbg_master_aw_burst[0]
port 791 nsew signal output
rlabel metal2 s 233146 359200 233202 360000 6 dbg_master_aw_burst[1]
port 792 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 dbg_master_aw_cache[0]
port 793 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 dbg_master_aw_cache[1]
port 794 nsew signal output
rlabel metal2 s 134614 359200 134670 360000 6 dbg_master_aw_cache[2]
port 795 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 dbg_master_aw_cache[3]
port 796 nsew signal output
rlabel metal3 s 0 206728 800 206848 6 dbg_master_aw_id[0]
port 797 nsew signal output
rlabel metal3 s 279200 286968 280000 287088 6 dbg_master_aw_id[1]
port 798 nsew signal output
rlabel metal3 s 0 246848 800 246968 6 dbg_master_aw_id[2]
port 799 nsew signal output
rlabel metal3 s 0 297168 800 297288 6 dbg_master_aw_id[3]
port 800 nsew signal output
rlabel metal2 s 226062 359200 226118 360000 6 dbg_master_aw_id[4]
port 801 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 dbg_master_aw_id[5]
port 802 nsew signal output
rlabel metal2 s 92754 359200 92810 360000 6 dbg_master_aw_id[6]
port 803 nsew signal output
rlabel metal3 s 0 240048 800 240168 6 dbg_master_aw_id[7]
port 804 nsew signal output
rlabel metal3 s 279200 207408 280000 207528 6 dbg_master_aw_id[8]
port 805 nsew signal output
rlabel metal3 s 0 210808 800 210928 6 dbg_master_aw_id[9]
port 806 nsew signal output
rlabel metal3 s 279200 174768 280000 174888 6 dbg_master_aw_len[0]
port 807 nsew signal output
rlabel metal3 s 0 305328 800 305448 6 dbg_master_aw_len[1]
port 808 nsew signal output
rlabel metal3 s 279200 159128 280000 159248 6 dbg_master_aw_len[2]
port 809 nsew signal output
rlabel metal2 s 101770 359200 101826 360000 6 dbg_master_aw_len[3]
port 810 nsew signal output
rlabel metal2 s 59910 359200 59966 360000 6 dbg_master_aw_len[4]
port 811 nsew signal output
rlabel metal2 s 273074 0 273130 800 6 dbg_master_aw_len[5]
port 812 nsew signal output
rlabel metal2 s 197082 359200 197138 360000 6 dbg_master_aw_len[6]
port 813 nsew signal output
rlabel metal2 s 245382 359200 245438 360000 6 dbg_master_aw_len[7]
port 814 nsew signal output
rlabel metal2 s 25134 359200 25190 360000 6 dbg_master_aw_lock
port 815 nsew signal output
rlabel metal2 s 256974 359200 257030 360000 6 dbg_master_aw_prot[0]
port 816 nsew signal output
rlabel metal2 s 38658 359200 38714 360000 6 dbg_master_aw_prot[1]
port 817 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 dbg_master_aw_prot[2]
port 818 nsew signal output
rlabel metal2 s 189998 359200 190054 360000 6 dbg_master_aw_qos[0]
port 819 nsew signal output
rlabel metal3 s 279200 268608 280000 268728 6 dbg_master_aw_qos[1]
port 820 nsew signal output
rlabel metal2 s 188066 359200 188122 360000 6 dbg_master_aw_qos[2]
port 821 nsew signal output
rlabel metal2 s 46386 359200 46442 360000 6 dbg_master_aw_qos[3]
port 822 nsew signal output
rlabel metal2 s 175830 359200 175886 360000 6 dbg_master_aw_ready
port 823 nsew signal input
rlabel metal3 s 279200 53728 280000 53848 6 dbg_master_aw_region[0]
port 824 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 dbg_master_aw_region[1]
port 825 nsew signal output
rlabel metal3 s 279200 191088 280000 191208 6 dbg_master_aw_region[2]
port 826 nsew signal output
rlabel metal3 s 279200 6808 280000 6928 6 dbg_master_aw_region[3]
port 827 nsew signal output
rlabel metal2 s 197726 359200 197782 360000 6 dbg_master_aw_size[0]
port 828 nsew signal output
rlabel metal3 s 279200 150288 280000 150408 6 dbg_master_aw_size[1]
port 829 nsew signal output
rlabel metal3 s 0 246168 800 246288 6 dbg_master_aw_size[2]
port 830 nsew signal output
rlabel metal3 s 0 324368 800 324488 6 dbg_master_aw_user[-1]
port 831 nsew signal output
rlabel metal3 s 0 358368 800 358488 6 dbg_master_aw_user[0]
port 832 nsew signal output
rlabel metal2 s 260194 359200 260250 360000 6 dbg_master_aw_valid
port 833 nsew signal output
rlabel metal2 s 200302 359200 200358 360000 6 dbg_master_b_id[0]
port 834 nsew signal input
rlabel metal3 s 279200 279488 280000 279608 6 dbg_master_b_id[1]
port 835 nsew signal input
rlabel metal3 s 279200 305328 280000 305448 6 dbg_master_b_id[2]
port 836 nsew signal input
rlabel metal2 s 122378 359200 122434 360000 6 dbg_master_b_id[3]
port 837 nsew signal input
rlabel metal3 s 0 350208 800 350328 6 dbg_master_b_id[4]
port 838 nsew signal input
rlabel metal3 s 279200 265208 280000 265328 6 dbg_master_b_id[5]
port 839 nsew signal input
rlabel metal2 s 199014 359200 199070 360000 6 dbg_master_b_id[6]
port 840 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 dbg_master_b_id[7]
port 841 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 dbg_master_b_id[8]
port 842 nsew signal input
rlabel metal3 s 279200 76168 280000 76288 6 dbg_master_b_id[9]
port 843 nsew signal input
rlabel metal3 s 0 278808 800 278928 6 dbg_master_b_ready
port 844 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 dbg_master_b_resp[0]
port 845 nsew signal input
rlabel metal2 s 168746 359200 168802 360000 6 dbg_master_b_resp[1]
port 846 nsew signal input
rlabel metal2 s 209962 359200 210018 360000 6 dbg_master_b_user[-1]
port 847 nsew signal input
rlabel metal2 s 190642 359200 190698 360000 6 dbg_master_b_user[0]
port 848 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 dbg_master_b_valid
port 849 nsew signal input
rlabel metal3 s 279200 354288 280000 354408 6 dbg_master_r_data[0]
port 850 nsew signal input
rlabel metal3 s 279200 280848 280000 280968 6 dbg_master_r_data[10]
port 851 nsew signal input
rlabel metal3 s 0 334568 800 334688 6 dbg_master_r_data[11]
port 852 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 dbg_master_r_data[12]
port 853 nsew signal input
rlabel metal3 s 0 145528 800 145648 6 dbg_master_r_data[13]
port 854 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 dbg_master_r_data[14]
port 855 nsew signal input
rlabel metal3 s 279200 159808 280000 159928 6 dbg_master_r_data[15]
port 856 nsew signal input
rlabel metal2 s 262770 0 262826 800 6 dbg_master_r_data[16]
port 857 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 dbg_master_r_data[17]
port 858 nsew signal input
rlabel metal3 s 279200 251608 280000 251728 6 dbg_master_r_data[18]
port 859 nsew signal input
rlabel metal2 s 106922 359200 106978 360000 6 dbg_master_r_data[19]
port 860 nsew signal input
rlabel metal3 s 279200 271328 280000 271448 6 dbg_master_r_data[1]
port 861 nsew signal input
rlabel metal3 s 279200 108128 280000 108248 6 dbg_master_r_data[20]
port 862 nsew signal input
rlabel metal2 s 51538 359200 51594 360000 6 dbg_master_r_data[21]
port 863 nsew signal input
rlabel metal2 s 45742 359200 45798 360000 6 dbg_master_r_data[22]
port 864 nsew signal input
rlabel metal2 s 128818 359200 128874 360000 6 dbg_master_r_data[23]
port 865 nsew signal input
rlabel metal2 s 138478 359200 138534 360000 6 dbg_master_r_data[24]
port 866 nsew signal input
rlabel metal2 s 263414 359200 263470 360000 6 dbg_master_r_data[25]
port 867 nsew signal input
rlabel metal2 s 120446 359200 120502 360000 6 dbg_master_r_data[26]
port 868 nsew signal input
rlabel metal3 s 279200 170008 280000 170128 6 dbg_master_r_data[27]
port 869 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 dbg_master_r_data[28]
port 870 nsew signal input
rlabel metal3 s 279200 65288 280000 65408 6 dbg_master_r_data[29]
port 871 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 dbg_master_r_data[2]
port 872 nsew signal input
rlabel metal2 s 123666 359200 123722 360000 6 dbg_master_r_data[30]
port 873 nsew signal input
rlabel metal3 s 0 184288 800 184408 6 dbg_master_r_data[31]
port 874 nsew signal input
rlabel metal2 s 244738 359200 244794 360000 6 dbg_master_r_data[32]
port 875 nsew signal input
rlabel metal2 s 117870 359200 117926 360000 6 dbg_master_r_data[33]
port 876 nsew signal input
rlabel metal2 s 246026 359200 246082 360000 6 dbg_master_r_data[34]
port 877 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 dbg_master_r_data[35]
port 878 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 dbg_master_r_data[36]
port 879 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 dbg_master_r_data[37]
port 880 nsew signal input
rlabel metal2 s 63130 359200 63186 360000 6 dbg_master_r_data[38]
port 881 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 dbg_master_r_data[39]
port 882 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 dbg_master_r_data[3]
port 883 nsew signal input
rlabel metal2 s 61198 359200 61254 360000 6 dbg_master_r_data[40]
port 884 nsew signal input
rlabel metal2 s 221554 359200 221610 360000 6 dbg_master_r_data[41]
port 885 nsew signal input
rlabel metal3 s 279200 236648 280000 236768 6 dbg_master_r_data[42]
port 886 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 dbg_master_r_data[43]
port 887 nsew signal input
rlabel metal3 s 0 330488 800 330608 6 dbg_master_r_data[44]
port 888 nsew signal input
rlabel metal2 s 73434 359200 73490 360000 6 dbg_master_r_data[45]
port 889 nsew signal input
rlabel metal3 s 279200 158448 280000 158568 6 dbg_master_r_data[46]
port 890 nsew signal input
rlabel metal2 s 237654 359200 237710 360000 6 dbg_master_r_data[47]
port 891 nsew signal input
rlabel metal2 s 111430 359200 111486 360000 6 dbg_master_r_data[48]
port 892 nsew signal input
rlabel metal2 s 70858 359200 70914 360000 6 dbg_master_r_data[49]
port 893 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 dbg_master_r_data[4]
port 894 nsew signal input
rlabel metal3 s 0 357688 800 357808 6 dbg_master_r_data[50]
port 895 nsew signal input
rlabel metal3 s 279200 8848 280000 8968 6 dbg_master_r_data[51]
port 896 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 dbg_master_r_data[52]
port 897 nsew signal input
rlabel metal3 s 279200 135328 280000 135448 6 dbg_master_r_data[53]
port 898 nsew signal input
rlabel metal3 s 0 172728 800 172848 6 dbg_master_r_data[54]
port 899 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 dbg_master_r_data[55]
port 900 nsew signal input
rlabel metal3 s 279200 34008 280000 34128 6 dbg_master_r_data[56]
port 901 nsew signal input
rlabel metal3 s 279200 355648 280000 355768 6 dbg_master_r_data[57]
port 902 nsew signal input
rlabel metal2 s 81806 359200 81862 360000 6 dbg_master_r_data[58]
port 903 nsew signal input
rlabel metal3 s 279200 356328 280000 356448 6 dbg_master_r_data[59]
port 904 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 dbg_master_r_data[5]
port 905 nsew signal input
rlabel metal3 s 0 357008 800 357128 6 dbg_master_r_data[60]
port 906 nsew signal input
rlabel metal2 s 230570 0 230626 800 6 dbg_master_r_data[61]
port 907 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 dbg_master_r_data[62]
port 908 nsew signal input
rlabel metal3 s 279200 289688 280000 289808 6 dbg_master_r_data[63]
port 909 nsew signal input
rlabel metal3 s 279200 329808 280000 329928 6 dbg_master_r_data[6]
port 910 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 dbg_master_r_data[7]
port 911 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 dbg_master_r_data[8]
port 912 nsew signal input
rlabel metal2 s 140410 359200 140466 360000 6 dbg_master_r_data[9]
port 913 nsew signal input
rlabel metal2 s 255042 0 255098 800 6 dbg_master_r_id[0]
port 914 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 dbg_master_r_id[1]
port 915 nsew signal input
rlabel metal3 s 0 257728 800 257848 6 dbg_master_r_id[2]
port 916 nsew signal input
rlabel metal3 s 0 255008 800 255128 6 dbg_master_r_id[3]
port 917 nsew signal input
rlabel metal2 s 210606 0 210662 800 6 dbg_master_r_id[4]
port 918 nsew signal input
rlabel metal2 s 257618 0 257674 800 6 dbg_master_r_id[5]
port 919 nsew signal input
rlabel metal3 s 279200 281528 280000 281648 6 dbg_master_r_id[6]
port 920 nsew signal input
rlabel metal3 s 279200 51688 280000 51808 6 dbg_master_r_id[7]
port 921 nsew signal input
rlabel metal3 s 0 274048 800 274168 6 dbg_master_r_id[8]
port 922 nsew signal input
rlabel metal3 s 279200 78888 280000 79008 6 dbg_master_r_id[9]
port 923 nsew signal input
rlabel metal3 s 279200 337288 280000 337408 6 dbg_master_r_last
port 924 nsew signal input
rlabel metal2 s 251178 0 251234 800 6 dbg_master_r_ready
port 925 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 dbg_master_r_resp[0]
port 926 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 dbg_master_r_resp[1]
port 927 nsew signal input
rlabel metal3 s 279200 235968 280000 236088 6 dbg_master_r_user[-1]
port 928 nsew signal input
rlabel metal3 s 279200 226448 280000 226568 6 dbg_master_r_user[0]
port 929 nsew signal input
rlabel metal3 s 0 208768 800 208888 6 dbg_master_r_valid
port 930 nsew signal input
rlabel metal3 s 279200 184288 280000 184408 6 dbg_master_w_data[0]
port 931 nsew signal output
rlabel metal3 s 0 189728 800 189848 6 dbg_master_w_data[10]
port 932 nsew signal output
rlabel metal2 s 159730 0 159786 800 6 dbg_master_w_data[11]
port 933 nsew signal output
rlabel metal3 s 0 146208 800 146328 6 dbg_master_w_data[12]
port 934 nsew signal output
rlabel metal3 s 279200 103368 280000 103488 6 dbg_master_w_data[13]
port 935 nsew signal output
rlabel metal2 s 274362 359200 274418 360000 6 dbg_master_w_data[14]
port 936 nsew signal output
rlabel metal2 s 180982 359200 181038 360000 6 dbg_master_w_data[15]
port 937 nsew signal output
rlabel metal3 s 0 316208 800 316328 6 dbg_master_w_data[16]
port 938 nsew signal output
rlabel metal2 s 220266 359200 220322 360000 6 dbg_master_w_data[17]
port 939 nsew signal output
rlabel metal3 s 0 271328 800 271448 6 dbg_master_w_data[18]
port 940 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 dbg_master_w_data[19]
port 941 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 dbg_master_w_data[1]
port 942 nsew signal output
rlabel metal3 s 0 337968 800 338088 6 dbg_master_w_data[20]
port 943 nsew signal output
rlabel metal2 s 279514 0 279570 800 6 dbg_master_w_data[21]
port 944 nsew signal output
rlabel metal3 s 279200 229168 280000 229288 6 dbg_master_w_data[22]
port 945 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 dbg_master_w_data[23]
port 946 nsew signal output
rlabel metal2 s 181626 359200 181682 360000 6 dbg_master_w_data[24]
port 947 nsew signal output
rlabel metal3 s 0 311448 800 311568 6 dbg_master_w_data[25]
port 948 nsew signal output
rlabel metal3 s 279200 113568 280000 113688 6 dbg_master_w_data[26]
port 949 nsew signal output
rlabel metal2 s 95330 359200 95386 360000 6 dbg_master_w_data[27]
port 950 nsew signal output
rlabel metal3 s 0 188368 800 188488 6 dbg_master_w_data[28]
port 951 nsew signal output
rlabel metal2 s 135258 359200 135314 360000 6 dbg_master_w_data[29]
port 952 nsew signal output
rlabel metal3 s 279200 100648 280000 100768 6 dbg_master_w_data[2]
port 953 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 dbg_master_w_data[30]
port 954 nsew signal output
rlabel metal3 s 0 325728 800 325848 6 dbg_master_w_data[31]
port 955 nsew signal output
rlabel metal3 s 279200 287648 280000 287768 6 dbg_master_w_data[32]
port 956 nsew signal output
rlabel metal3 s 0 318928 800 319048 6 dbg_master_w_data[33]
port 957 nsew signal output
rlabel metal2 s 15474 359200 15530 360000 6 dbg_master_w_data[34]
port 958 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 dbg_master_w_data[35]
port 959 nsew signal output
rlabel metal3 s 279200 344088 280000 344208 6 dbg_master_w_data[36]
port 960 nsew signal output
rlabel metal2 s 253110 359200 253166 360000 6 dbg_master_w_data[37]
port 961 nsew signal output
rlabel metal3 s 279200 163888 280000 164008 6 dbg_master_w_data[38]
port 962 nsew signal output
rlabel metal3 s 0 240728 800 240848 6 dbg_master_w_data[39]
port 963 nsew signal output
rlabel metal3 s 0 150288 800 150408 6 dbg_master_w_data[3]
port 964 nsew signal output
rlabel metal3 s 279200 211488 280000 211608 6 dbg_master_w_data[40]
port 965 nsew signal output
rlabel metal3 s 0 238688 800 238808 6 dbg_master_w_data[41]
port 966 nsew signal output
rlabel metal3 s 0 283568 800 283688 6 dbg_master_w_data[42]
port 967 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 dbg_master_w_data[43]
port 968 nsew signal output
rlabel metal2 s 32862 359200 32918 360000 6 dbg_master_w_data[44]
port 969 nsew signal output
rlabel metal3 s 279200 304648 280000 304768 6 dbg_master_w_data[45]
port 970 nsew signal output
rlabel metal2 s 237654 0 237710 800 6 dbg_master_w_data[46]
port 971 nsew signal output
rlabel metal3 s 0 260448 800 260568 6 dbg_master_w_data[47]
port 972 nsew signal output
rlabel metal3 s 279200 208088 280000 208208 6 dbg_master_w_data[48]
port 973 nsew signal output
rlabel metal2 s 106278 359200 106334 360000 6 dbg_master_w_data[49]
port 974 nsew signal output
rlabel metal2 s 269854 0 269910 800 6 dbg_master_w_data[4]
port 975 nsew signal output
rlabel metal3 s 0 342728 800 342848 6 dbg_master_w_data[50]
port 976 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 dbg_master_w_data[51]
port 977 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 dbg_master_w_data[52]
port 978 nsew signal output
rlabel metal3 s 0 348168 800 348288 6 dbg_master_w_data[53]
port 979 nsew signal output
rlabel metal2 s 68282 359200 68338 360000 6 dbg_master_w_data[54]
port 980 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 dbg_master_w_data[55]
port 981 nsew signal output
rlabel metal2 s 18694 359200 18750 360000 6 dbg_master_w_data[56]
port 982 nsew signal output
rlabel metal3 s 0 149608 800 149728 6 dbg_master_w_data[57]
port 983 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 dbg_master_w_data[58]
port 984 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 dbg_master_w_data[59]
port 985 nsew signal output
rlabel metal3 s 0 157768 800 157888 6 dbg_master_w_data[5]
port 986 nsew signal output
rlabel metal3 s 0 159128 800 159248 6 dbg_master_w_data[60]
port 987 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 dbg_master_w_data[61]
port 988 nsew signal output
rlabel metal2 s 193862 0 193918 800 6 dbg_master_w_data[62]
port 989 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 dbg_master_w_data[63]
port 990 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 dbg_master_w_data[6]
port 991 nsew signal output
rlabel metal2 s 254398 359200 254454 360000 6 dbg_master_w_data[7]
port 992 nsew signal output
rlabel metal3 s 0 688 800 808 6 dbg_master_w_data[8]
port 993 nsew signal output
rlabel metal2 s 213826 359200 213882 360000 6 dbg_master_w_data[9]
port 994 nsew signal output
rlabel metal3 s 0 162528 800 162648 6 dbg_master_w_last
port 995 nsew signal output
rlabel metal2 s 276294 0 276350 800 6 dbg_master_w_ready
port 996 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 dbg_master_w_strb[0]
port 997 nsew signal output
rlabel metal2 s 84382 359200 84438 360000 6 dbg_master_w_strb[1]
port 998 nsew signal output
rlabel metal3 s 279200 326408 280000 326528 6 dbg_master_w_strb[2]
port 999 nsew signal output
rlabel metal3 s 0 268608 800 268728 6 dbg_master_w_strb[3]
port 1000 nsew signal output
rlabel metal3 s 279200 320968 280000 321088 6 dbg_master_w_strb[4]
port 1001 nsew signal output
rlabel metal3 s 279200 53048 280000 53168 6 dbg_master_w_strb[5]
port 1002 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 dbg_master_w_strb[6]
port 1003 nsew signal output
rlabel metal3 s 279200 194488 280000 194608 6 dbg_master_w_strb[7]
port 1004 nsew signal output
rlabel metal3 s 279200 142128 280000 142248 6 dbg_master_w_user[-1]
port 1005 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 dbg_master_w_user[0]
port 1006 nsew signal output
rlabel metal2 s 14186 359200 14242 360000 6 dbg_master_w_valid
port 1007 nsew signal output
rlabel metal3 s 279200 144848 280000 144968 6 debug_addr[0]
port 1008 nsew signal input
rlabel metal2 s 16762 359200 16818 360000 6 debug_addr[10]
port 1009 nsew signal input
rlabel metal3 s 0 267928 800 268048 6 debug_addr[11]
port 1010 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 debug_addr[12]
port 1011 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 debug_addr[13]
port 1012 nsew signal input
rlabel metal2 s 269210 359200 269266 360000 6 debug_addr[14]
port 1013 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 debug_addr[1]
port 1014 nsew signal input
rlabel metal3 s 0 216928 800 217048 6 debug_addr[2]
port 1015 nsew signal input
rlabel metal3 s 279200 199928 280000 200048 6 debug_addr[3]
port 1016 nsew signal input
rlabel metal3 s 0 293088 800 293208 6 debug_addr[4]
port 1017 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 debug_addr[5]
port 1018 nsew signal input
rlabel metal3 s 279200 180888 280000 181008 6 debug_addr[6]
port 1019 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 debug_addr[7]
port 1020 nsew signal input
rlabel metal3 s 279200 234608 280000 234728 6 debug_addr[8]
port 1021 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 debug_addr[9]
port 1022 nsew signal input
rlabel metal3 s 279200 123088 280000 123208 6 debug_gnt
port 1023 nsew signal output
rlabel metal2 s 269854 359200 269910 360000 6 debug_rdata[0]
port 1024 nsew signal output
rlabel metal3 s 279200 93848 280000 93968 6 debug_rdata[10]
port 1025 nsew signal output
rlabel metal3 s 0 299208 800 299328 6 debug_rdata[11]
port 1026 nsew signal output
rlabel metal2 s 211250 359200 211306 360000 6 debug_rdata[12]
port 1027 nsew signal output
rlabel metal3 s 279200 192448 280000 192568 6 debug_rdata[13]
port 1028 nsew signal output
rlabel metal2 s 137190 359200 137246 360000 6 debug_rdata[14]
port 1029 nsew signal output
rlabel metal2 s 276938 0 276994 800 6 debug_rdata[15]
port 1030 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 debug_rdata[16]
port 1031 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 debug_rdata[17]
port 1032 nsew signal output
rlabel metal3 s 0 161168 800 161288 6 debug_rdata[18]
port 1033 nsew signal output
rlabel metal3 s 279200 202648 280000 202768 6 debug_rdata[19]
port 1034 nsew signal output
rlabel metal2 s 193862 359200 193918 360000 6 debug_rdata[1]
port 1035 nsew signal output
rlabel metal3 s 279200 189048 280000 189168 6 debug_rdata[20]
port 1036 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 debug_rdata[21]
port 1037 nsew signal output
rlabel metal3 s 279200 17688 280000 17808 6 debug_rdata[22]
port 1038 nsew signal output
rlabel metal3 s 279200 216928 280000 217048 6 debug_rdata[23]
port 1039 nsew signal output
rlabel metal3 s 279200 46928 280000 47048 6 debug_rdata[24]
port 1040 nsew signal output
rlabel metal3 s 279200 71408 280000 71528 6 debug_rdata[25]
port 1041 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 debug_rdata[26]
port 1042 nsew signal output
rlabel metal2 s 259550 0 259606 800 6 debug_rdata[27]
port 1043 nsew signal output
rlabel metal3 s 279200 79568 280000 79688 6 debug_rdata[28]
port 1044 nsew signal output
rlabel metal2 s 28998 359200 29054 360000 6 debug_rdata[29]
port 1045 nsew signal output
rlabel metal3 s 279200 94528 280000 94648 6 debug_rdata[2]
port 1046 nsew signal output
rlabel metal3 s 0 310768 800 310888 6 debug_rdata[30]
port 1047 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 debug_rdata[31]
port 1048 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 debug_rdata[3]
port 1049 nsew signal output
rlabel metal2 s 48962 359200 49018 360000 6 debug_rdata[4]
port 1050 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 debug_rdata[5]
port 1051 nsew signal output
rlabel metal3 s 279200 266568 280000 266688 6 debug_rdata[6]
port 1052 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 debug_rdata[7]
port 1053 nsew signal output
rlabel metal2 s 252466 359200 252522 360000 6 debug_rdata[8]
port 1054 nsew signal output
rlabel metal2 s 235722 0 235778 800 6 debug_rdata[9]
port 1055 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 debug_req
port 1056 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 debug_rvalid
port 1057 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 debug_wdata[0]
port 1058 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 debug_wdata[10]
port 1059 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 debug_wdata[11]
port 1060 nsew signal input
rlabel metal2 s 260194 0 260250 800 6 debug_wdata[12]
port 1061 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 debug_wdata[13]
port 1062 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 debug_wdata[14]
port 1063 nsew signal input
rlabel metal2 s 1950 359200 2006 360000 6 debug_wdata[15]
port 1064 nsew signal input
rlabel metal2 s 36726 359200 36782 360000 6 debug_wdata[16]
port 1065 nsew signal input
rlabel metal2 s 70214 359200 70270 360000 6 debug_wdata[17]
port 1066 nsew signal input
rlabel metal3 s 279200 162528 280000 162648 6 debug_wdata[18]
port 1067 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 debug_wdata[19]
port 1068 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 debug_wdata[1]
port 1069 nsew signal input
rlabel metal3 s 0 194488 800 194608 6 debug_wdata[20]
port 1070 nsew signal input
rlabel metal3 s 279200 297848 280000 297968 6 debug_wdata[21]
port 1071 nsew signal input
rlabel metal3 s 279200 201968 280000 202088 6 debug_wdata[22]
port 1072 nsew signal input
rlabel metal3 s 279200 59168 280000 59288 6 debug_wdata[23]
port 1073 nsew signal input
rlabel metal3 s 279200 156408 280000 156528 6 debug_wdata[24]
port 1074 nsew signal input
rlabel metal3 s 279200 240728 280000 240848 6 debug_wdata[25]
port 1075 nsew signal input
rlabel metal3 s 279200 306688 280000 306808 6 debug_wdata[26]
port 1076 nsew signal input
rlabel metal3 s 279200 126488 280000 126608 6 debug_wdata[27]
port 1077 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 debug_wdata[28]
port 1078 nsew signal input
rlabel metal3 s 279200 227128 280000 227248 6 debug_wdata[29]
port 1079 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 debug_wdata[2]
port 1080 nsew signal input
rlabel metal2 s 173898 359200 173954 360000 6 debug_wdata[30]
port 1081 nsew signal input
rlabel metal3 s 279200 246848 280000 246968 6 debug_wdata[31]
port 1082 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 debug_wdata[3]
port 1083 nsew signal input
rlabel metal3 s 279200 292408 280000 292528 6 debug_wdata[4]
port 1084 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 debug_wdata[5]
port 1085 nsew signal input
rlabel metal3 s 279200 157088 280000 157208 6 debug_wdata[6]
port 1086 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 debug_wdata[7]
port 1087 nsew signal input
rlabel metal2 s 195794 0 195850 800 6 debug_wdata[8]
port 1088 nsew signal input
rlabel metal3 s 279200 69368 280000 69488 6 debug_wdata[9]
port 1089 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 debug_we
port 1090 nsew signal input
rlabel metal2 s 182914 359200 182970 360000 6 fetch_enable_i
port 1091 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 instr_slave_ar_addr[0]
port 1092 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 instr_slave_ar_addr[10]
port 1093 nsew signal input
rlabel metal3 s 0 252968 800 253088 6 instr_slave_ar_addr[11]
port 1094 nsew signal input
rlabel metal3 s 279200 276088 280000 276208 6 instr_slave_ar_addr[12]
port 1095 nsew signal input
rlabel metal3 s 279200 283568 280000 283688 6 instr_slave_ar_addr[13]
port 1096 nsew signal input
rlabel metal3 s 279200 60528 280000 60648 6 instr_slave_ar_addr[14]
port 1097 nsew signal input
rlabel metal2 s 240874 359200 240930 360000 6 instr_slave_ar_addr[15]
port 1098 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 instr_slave_ar_addr[16]
port 1099 nsew signal input
rlabel metal2 s 139122 359200 139178 360000 6 instr_slave_ar_addr[17]
port 1100 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 instr_slave_ar_addr[18]
port 1101 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 instr_slave_ar_addr[19]
port 1102 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 instr_slave_ar_addr[1]
port 1103 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 instr_slave_ar_addr[20]
port 1104 nsew signal input
rlabel metal3 s 279200 329128 280000 329248 6 instr_slave_ar_addr[21]
port 1105 nsew signal input
rlabel metal3 s 279200 72768 280000 72888 6 instr_slave_ar_addr[22]
port 1106 nsew signal input
rlabel metal2 s 27066 359200 27122 360000 6 instr_slave_ar_addr[23]
port 1107 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 instr_slave_ar_addr[24]
port 1108 nsew signal input
rlabel metal3 s 0 350888 800 351008 6 instr_slave_ar_addr[25]
port 1109 nsew signal input
rlabel metal3 s 0 310088 800 310208 6 instr_slave_ar_addr[26]
port 1110 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 instr_slave_ar_addr[27]
port 1111 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 instr_slave_ar_addr[28]
port 1112 nsew signal input
rlabel metal3 s 279200 308048 280000 308168 6 instr_slave_ar_addr[29]
port 1113 nsew signal input
rlabel metal3 s 279200 140768 280000 140888 6 instr_slave_ar_addr[2]
port 1114 nsew signal input
rlabel metal2 s 123022 359200 123078 360000 6 instr_slave_ar_addr[30]
port 1115 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 instr_slave_ar_addr[31]
port 1116 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 instr_slave_ar_addr[3]
port 1117 nsew signal input
rlabel metal3 s 279200 320288 280000 320408 6 instr_slave_ar_addr[4]
port 1118 nsew signal input
rlabel metal3 s 0 275408 800 275528 6 instr_slave_ar_addr[5]
port 1119 nsew signal input
rlabel metal3 s 279200 246168 280000 246288 6 instr_slave_ar_addr[6]
port 1120 nsew signal input
rlabel metal3 s 279200 299888 280000 300008 6 instr_slave_ar_addr[7]
port 1121 nsew signal input
rlabel metal3 s 279200 164568 280000 164688 6 instr_slave_ar_addr[8]
port 1122 nsew signal input
rlabel metal3 s 279200 54408 280000 54528 6 instr_slave_ar_addr[9]
port 1123 nsew signal input
rlabel metal3 s 279200 157768 280000 157888 6 instr_slave_ar_burst[0]
port 1124 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 instr_slave_ar_burst[1]
port 1125 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 instr_slave_ar_cache[0]
port 1126 nsew signal input
rlabel metal3 s 0 174088 800 174208 6 instr_slave_ar_cache[1]
port 1127 nsew signal input
rlabel metal2 s 10966 359200 11022 360000 6 instr_slave_ar_cache[2]
port 1128 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 instr_slave_ar_cache[3]
port 1129 nsew signal input
rlabel metal3 s 279200 238688 280000 238808 6 instr_slave_ar_id[0]
port 1130 nsew signal input
rlabel metal2 s 115938 359200 115994 360000 6 instr_slave_ar_id[1]
port 1131 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 instr_slave_ar_id[2]
port 1132 nsew signal input
rlabel metal3 s 0 228488 800 228608 6 instr_slave_ar_id[3]
port 1133 nsew signal input
rlabel metal2 s 272430 359200 272486 360000 6 instr_slave_ar_id[4]
port 1134 nsew signal input
rlabel metal2 s 79874 359200 79930 360000 6 instr_slave_ar_id[5]
port 1135 nsew signal input
rlabel metal3 s 279200 155048 280000 155168 6 instr_slave_ar_id[6]
port 1136 nsew signal input
rlabel metal3 s 0 317568 800 317688 6 instr_slave_ar_id[7]
port 1137 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 instr_slave_ar_id[8]
port 1138 nsew signal input
rlabel metal3 s 0 197888 800 198008 6 instr_slave_ar_id[9]
port 1139 nsew signal input
rlabel metal3 s 279200 15648 280000 15768 6 instr_slave_ar_len[0]
port 1140 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 instr_slave_ar_len[1]
port 1141 nsew signal input
rlabel metal3 s 0 259088 800 259208 6 instr_slave_ar_len[2]
port 1142 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 instr_slave_ar_len[3]
port 1143 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 instr_slave_ar_len[4]
port 1144 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 instr_slave_ar_len[5]
port 1145 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 instr_slave_ar_len[6]
port 1146 nsew signal input
rlabel metal2 s 191286 359200 191342 360000 6 instr_slave_ar_len[7]
port 1147 nsew signal input
rlabel metal3 s 279200 219648 280000 219768 6 instr_slave_ar_lock
port 1148 nsew signal input
rlabel metal2 s 208030 359200 208086 360000 6 instr_slave_ar_prot[0]
port 1149 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 instr_slave_ar_prot[1]
port 1150 nsew signal input
rlabel metal3 s 0 242768 800 242888 6 instr_slave_ar_prot[2]
port 1151 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 instr_slave_ar_qos[0]
port 1152 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 instr_slave_ar_qos[1]
port 1153 nsew signal input
rlabel metal3 s 0 284248 800 284368 6 instr_slave_ar_qos[2]
port 1154 nsew signal input
rlabel metal2 s 272430 0 272486 800 6 instr_slave_ar_qos[3]
port 1155 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 instr_slave_ar_ready
port 1156 nsew signal output
rlabel metal3 s 279200 294448 280000 294568 6 instr_slave_ar_region[0]
port 1157 nsew signal input
rlabel metal3 s 279200 212848 280000 212968 6 instr_slave_ar_region[1]
port 1158 nsew signal input
rlabel metal3 s 279200 90448 280000 90568 6 instr_slave_ar_region[2]
port 1159 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 instr_slave_ar_region[3]
port 1160 nsew signal input
rlabel metal3 s 279200 214888 280000 215008 6 instr_slave_ar_size[0]
port 1161 nsew signal input
rlabel metal3 s 0 167968 800 168088 6 instr_slave_ar_size[1]
port 1162 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 instr_slave_ar_size[2]
port 1163 nsew signal input
rlabel metal3 s 0 201968 800 202088 6 instr_slave_ar_user[-1]
port 1164 nsew signal input
rlabel metal2 s 158442 359200 158498 360000 6 instr_slave_ar_user[0]
port 1165 nsew signal input
rlabel metal3 s 0 308048 800 308168 6 instr_slave_ar_valid
port 1166 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 instr_slave_aw_addr[0]
port 1167 nsew signal input
rlabel metal2 s 232502 359200 232558 360000 6 instr_slave_aw_addr[10]
port 1168 nsew signal input
rlabel metal3 s 279200 55768 280000 55888 6 instr_slave_aw_addr[11]
port 1169 nsew signal input
rlabel metal3 s 279200 328448 280000 328568 6 instr_slave_aw_addr[12]
port 1170 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 instr_slave_aw_addr[13]
port 1171 nsew signal input
rlabel metal3 s 279200 282208 280000 282328 6 instr_slave_aw_addr[14]
port 1172 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 instr_slave_aw_addr[15]
port 1173 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 instr_slave_aw_addr[16]
port 1174 nsew signal input
rlabel metal3 s 279200 264528 280000 264648 6 instr_slave_aw_addr[17]
port 1175 nsew signal input
rlabel metal3 s 279200 151648 280000 151768 6 instr_slave_aw_addr[18]
port 1176 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 instr_slave_aw_addr[19]
port 1177 nsew signal input
rlabel metal3 s 279200 161848 280000 161968 6 instr_slave_aw_addr[1]
port 1178 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 instr_slave_aw_addr[20]
port 1179 nsew signal input
rlabel metal2 s 125598 359200 125654 360000 6 instr_slave_aw_addr[21]
port 1180 nsew signal input
rlabel metal3 s 279200 252968 280000 253088 6 instr_slave_aw_addr[22]
port 1181 nsew signal input
rlabel metal3 s 0 172048 800 172168 6 instr_slave_aw_addr[23]
port 1182 nsew signal input
rlabel metal2 s 217690 0 217746 800 6 instr_slave_aw_addr[24]
port 1183 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 instr_slave_aw_addr[25]
port 1184 nsew signal input
rlabel metal3 s 279200 81608 280000 81728 6 instr_slave_aw_addr[26]
port 1185 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 instr_slave_aw_addr[27]
port 1186 nsew signal input
rlabel metal3 s 0 286968 800 287088 6 instr_slave_aw_addr[28]
port 1187 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 instr_slave_aw_addr[29]
port 1188 nsew signal input
rlabel metal3 s 279200 203328 280000 203448 6 instr_slave_aw_addr[2]
port 1189 nsew signal input
rlabel metal3 s 279200 28568 280000 28688 6 instr_slave_aw_addr[30]
port 1190 nsew signal input
rlabel metal3 s 279200 345448 280000 345568 6 instr_slave_aw_addr[31]
port 1191 nsew signal input
rlabel metal3 s 279200 340008 280000 340128 6 instr_slave_aw_addr[3]
port 1192 nsew signal input
rlabel metal3 s 0 187688 800 187808 6 instr_slave_aw_addr[4]
port 1193 nsew signal input
rlabel metal3 s 279200 336608 280000 336728 6 instr_slave_aw_addr[5]
port 1194 nsew signal input
rlabel metal2 s 171322 359200 171378 360000 6 instr_slave_aw_addr[6]
port 1195 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 instr_slave_aw_addr[7]
port 1196 nsew signal input
rlabel metal2 s 23202 359200 23258 360000 6 instr_slave_aw_addr[8]
port 1197 nsew signal input
rlabel metal2 s 144274 359200 144330 360000 6 instr_slave_aw_addr[9]
port 1198 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 instr_slave_aw_burst[0]
port 1199 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 instr_slave_aw_burst[1]
port 1200 nsew signal input
rlabel metal3 s 0 259768 800 259888 6 instr_slave_aw_cache[0]
port 1201 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 instr_slave_aw_cache[1]
port 1202 nsew signal input
rlabel metal3 s 279200 31288 280000 31408 6 instr_slave_aw_cache[2]
port 1203 nsew signal input
rlabel metal3 s 0 256368 800 256488 6 instr_slave_aw_cache[3]
port 1204 nsew signal input
rlabel metal3 s 279200 318248 280000 318368 6 instr_slave_aw_id[0]
port 1205 nsew signal input
rlabel metal3 s 279200 267248 280000 267368 6 instr_slave_aw_id[1]
port 1206 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 instr_slave_aw_id[2]
port 1207 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 instr_slave_aw_id[3]
port 1208 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 instr_slave_aw_id[4]
port 1209 nsew signal input
rlabel metal3 s 279200 227808 280000 227928 6 instr_slave_aw_id[5]
port 1210 nsew signal input
rlabel metal2 s 90178 359200 90234 360000 6 instr_slave_aw_id[6]
port 1211 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 instr_slave_aw_id[7]
port 1212 nsew signal input
rlabel metal2 s 163594 359200 163650 360000 6 instr_slave_aw_id[8]
port 1213 nsew signal input
rlabel metal2 s 7746 359200 7802 360000 6 instr_slave_aw_id[9]
port 1214 nsew signal input
rlabel metal3 s 279200 68008 280000 68128 6 instr_slave_aw_len[0]
port 1215 nsew signal input
rlabel metal3 s 279200 218968 280000 219088 6 instr_slave_aw_len[1]
port 1216 nsew signal input
rlabel metal3 s 0 295128 800 295248 6 instr_slave_aw_len[2]
port 1217 nsew signal input
rlabel metal3 s 0 231888 800 232008 6 instr_slave_aw_len[3]
port 1218 nsew signal input
rlabel metal3 s 279200 153008 280000 153128 6 instr_slave_aw_len[4]
port 1219 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 instr_slave_aw_len[5]
port 1220 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 instr_slave_aw_len[6]
port 1221 nsew signal input
rlabel metal2 s 152646 359200 152702 360000 6 instr_slave_aw_len[7]
port 1222 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 instr_slave_aw_lock
port 1223 nsew signal input
rlabel metal3 s 0 185648 800 185768 6 instr_slave_aw_prot[0]
port 1224 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 instr_slave_aw_prot[1]
port 1225 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 instr_slave_aw_prot[2]
port 1226 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 instr_slave_aw_qos[0]
port 1227 nsew signal input
rlabel metal2 s 147494 359200 147550 360000 6 instr_slave_aw_qos[1]
port 1228 nsew signal input
rlabel metal2 s 34150 359200 34206 360000 6 instr_slave_aw_qos[2]
port 1229 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 instr_slave_aw_qos[3]
port 1230 nsew signal input
rlabel metal3 s 279200 239368 280000 239488 6 instr_slave_aw_ready
port 1231 nsew signal output
rlabel metal2 s 44454 359200 44510 360000 6 instr_slave_aw_region[0]
port 1232 nsew signal input
rlabel metal3 s 279200 221688 280000 221808 6 instr_slave_aw_region[1]
port 1233 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 instr_slave_aw_region[2]
port 1234 nsew signal input
rlabel metal3 s 279200 14288 280000 14408 6 instr_slave_aw_region[3]
port 1235 nsew signal input
rlabel metal2 s 75366 359200 75422 360000 6 instr_slave_aw_size[0]
port 1236 nsew signal input
rlabel metal3 s 0 303968 800 304088 6 instr_slave_aw_size[1]
port 1237 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 instr_slave_aw_size[2]
port 1238 nsew signal input
rlabel metal2 s 234434 359200 234490 360000 6 instr_slave_aw_user[-1]
port 1239 nsew signal input
rlabel metal3 s 279200 52368 280000 52488 6 instr_slave_aw_user[0]
port 1240 nsew signal input
rlabel metal2 s 112074 359200 112130 360000 6 instr_slave_aw_valid
port 1241 nsew signal input
rlabel metal2 s 83094 359200 83150 360000 6 instr_slave_b_id[0]
port 1242 nsew signal output
rlabel metal2 s 249890 0 249946 800 6 instr_slave_b_id[1]
port 1243 nsew signal output
rlabel metal3 s 0 309408 800 309528 6 instr_slave_b_id[2]
port 1244 nsew signal output
rlabel metal3 s 0 209448 800 209568 6 instr_slave_b_id[3]
port 1245 nsew signal output
rlabel metal2 s 57978 359200 58034 360000 6 instr_slave_b_id[4]
port 1246 nsew signal output
rlabel metal2 s 8390 359200 8446 360000 6 instr_slave_b_id[5]
port 1247 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 instr_slave_b_id[6]
port 1248 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 instr_slave_b_id[7]
port 1249 nsew signal output
rlabel metal3 s 279200 316888 280000 317008 6 instr_slave_b_id[8]
port 1250 nsew signal output
rlabel metal2 s 209318 359200 209374 360000 6 instr_slave_b_id[9]
port 1251 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 instr_slave_b_ready
port 1252 nsew signal input
rlabel metal3 s 0 319608 800 319728 6 instr_slave_b_resp[0]
port 1253 nsew signal output
rlabel metal2 s 253110 0 253166 800 6 instr_slave_b_resp[1]
port 1254 nsew signal output
rlabel metal3 s 279200 179528 280000 179648 6 instr_slave_b_user[-1]
port 1255 nsew signal output
rlabel metal2 s 247958 359200 248014 360000 6 instr_slave_b_user[0]
port 1256 nsew signal output
rlabel metal2 s 208030 0 208086 800 6 instr_slave_b_valid
port 1257 nsew signal output
rlabel metal3 s 0 204688 800 204808 6 instr_slave_r_data[0]
port 1258 nsew signal output
rlabel metal2 s 118514 359200 118570 360000 6 instr_slave_r_data[10]
port 1259 nsew signal output
rlabel metal3 s 279200 175448 280000 175568 6 instr_slave_r_data[11]
port 1260 nsew signal output
rlabel metal3 s 279200 344768 280000 344888 6 instr_slave_r_data[12]
port 1261 nsew signal output
rlabel metal3 s 279200 257728 280000 257848 6 instr_slave_r_data[13]
port 1262 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 instr_slave_r_data[14]
port 1263 nsew signal output
rlabel metal3 s 0 233928 800 234048 6 instr_slave_r_data[15]
port 1264 nsew signal output
rlabel metal3 s 279200 40128 280000 40248 6 instr_slave_r_data[16]
port 1265 nsew signal output
rlabel metal2 s 177118 359200 177174 360000 6 instr_slave_r_data[17]
port 1266 nsew signal output
rlabel metal3 s 279200 122408 280000 122528 6 instr_slave_r_data[18]
port 1267 nsew signal output
rlabel metal3 s 279200 312128 280000 312248 6 instr_slave_r_data[19]
port 1268 nsew signal output
rlabel metal2 s 74078 359200 74134 360000 6 instr_slave_r_data[1]
port 1269 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 instr_slave_r_data[20]
port 1270 nsew signal output
rlabel metal3 s 279200 174088 280000 174208 6 instr_slave_r_data[21]
port 1271 nsew signal output
rlabel metal3 s 279200 84328 280000 84448 6 instr_slave_r_data[22]
port 1272 nsew signal output
rlabel metal2 s 3882 359200 3938 360000 6 instr_slave_r_data[23]
port 1273 nsew signal output
rlabel metal2 s 9034 359200 9090 360000 6 instr_slave_r_data[24]
port 1274 nsew signal output
rlabel metal3 s 279200 275408 280000 275528 6 instr_slave_r_data[25]
port 1275 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 instr_slave_r_data[26]
port 1276 nsew signal output
rlabel metal2 s 229282 0 229338 800 6 instr_slave_r_data[27]
port 1277 nsew signal output
rlabel metal2 s 242806 0 242862 800 6 instr_slave_r_data[28]
port 1278 nsew signal output
rlabel metal3 s 279200 322328 280000 322448 6 instr_slave_r_data[29]
port 1279 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 instr_slave_r_data[2]
port 1280 nsew signal output
rlabel metal3 s 279200 198568 280000 198688 6 instr_slave_r_data[30]
port 1281 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 instr_slave_r_data[31]
port 1282 nsew signal output
rlabel metal3 s 279200 233248 280000 233368 6 instr_slave_r_data[32]
port 1283 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 instr_slave_r_data[33]
port 1284 nsew signal output
rlabel metal3 s 279200 4088 280000 4208 6 instr_slave_r_data[34]
port 1285 nsew signal output
rlabel metal3 s 279200 346128 280000 346248 6 instr_slave_r_data[35]
port 1286 nsew signal output
rlabel metal2 s 233790 359200 233846 360000 6 instr_slave_r_data[36]
port 1287 nsew signal output
rlabel metal2 s 114006 359200 114062 360000 6 instr_slave_r_data[37]
port 1288 nsew signal output
rlabel metal2 s 210606 359200 210662 360000 6 instr_slave_r_data[38]
port 1289 nsew signal output
rlabel metal3 s 0 236648 800 236768 6 instr_slave_r_data[39]
port 1290 nsew signal output
rlabel metal3 s 279200 63248 280000 63368 6 instr_slave_r_data[3]
port 1291 nsew signal output
rlabel metal2 s 207386 359200 207442 360000 6 instr_slave_r_data[40]
port 1292 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 instr_slave_r_data[41]
port 1293 nsew signal output
rlabel metal3 s 279200 23808 280000 23928 6 instr_slave_r_data[42]
port 1294 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 instr_slave_r_data[43]
port 1295 nsew signal output
rlabel metal2 s 220910 0 220966 800 6 instr_slave_r_data[44]
port 1296 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 instr_slave_r_data[45]
port 1297 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 instr_slave_r_data[46]
port 1298 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 instr_slave_r_data[47]
port 1299 nsew signal output
rlabel metal2 s 209318 0 209374 800 6 instr_slave_r_data[48]
port 1300 nsew signal output
rlabel metal3 s 0 204008 800 204128 6 instr_slave_r_data[49]
port 1301 nsew signal output
rlabel metal3 s 0 293768 800 293888 6 instr_slave_r_data[4]
port 1302 nsew signal output
rlabel metal3 s 279200 148248 280000 148368 6 instr_slave_r_data[50]
port 1303 nsew signal output
rlabel metal3 s 0 167288 800 167408 6 instr_slave_r_data[51]
port 1304 nsew signal output
rlabel metal3 s 279200 184968 280000 185088 6 instr_slave_r_data[52]
port 1305 nsew signal output
rlabel metal3 s 279200 248208 280000 248328 6 instr_slave_r_data[53]
port 1306 nsew signal output
rlabel metal3 s 279200 7488 280000 7608 6 instr_slave_r_data[54]
port 1307 nsew signal output
rlabel metal3 s 0 252288 800 252408 6 instr_slave_r_data[55]
port 1308 nsew signal output
rlabel metal2 s 266634 0 266690 800 6 instr_slave_r_data[56]
port 1309 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 instr_slave_r_data[57]
port 1310 nsew signal output
rlabel metal3 s 0 342048 800 342168 6 instr_slave_r_data[58]
port 1311 nsew signal output
rlabel metal2 s 275006 359200 275062 360000 6 instr_slave_r_data[59]
port 1312 nsew signal output
rlabel metal2 s 12898 359200 12954 360000 6 instr_slave_r_data[5]
port 1313 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 instr_slave_r_data[60]
port 1314 nsew signal output
rlabel metal3 s 279200 75488 280000 75608 6 instr_slave_r_data[61]
port 1315 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 instr_slave_r_data[62]
port 1316 nsew signal output
rlabel metal3 s 279200 284928 280000 285048 6 instr_slave_r_data[63]
port 1317 nsew signal output
rlabel metal3 s 279200 311448 280000 311568 6 instr_slave_r_data[6]
port 1318 nsew signal output
rlabel metal2 s 265990 359200 266046 360000 6 instr_slave_r_data[7]
port 1319 nsew signal output
rlabel metal2 s 47030 359200 47086 360000 6 instr_slave_r_data[8]
port 1320 nsew signal output
rlabel metal2 s 154578 359200 154634 360000 6 instr_slave_r_data[9]
port 1321 nsew signal output
rlabel metal3 s 0 218968 800 219088 6 instr_slave_r_id[0]
port 1322 nsew signal output
rlabel metal2 s 10322 359200 10378 360000 6 instr_slave_r_id[1]
port 1323 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 instr_slave_r_id[2]
port 1324 nsew signal output
rlabel metal2 s 89534 359200 89590 360000 6 instr_slave_r_id[3]
port 1325 nsew signal output
rlabel metal3 s 279200 350888 280000 351008 6 instr_slave_r_id[4]
port 1326 nsew signal output
rlabel metal2 s 52826 359200 52882 360000 6 instr_slave_r_id[5]
port 1327 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 instr_slave_r_id[6]
port 1328 nsew signal output
rlabel metal3 s 279200 112208 280000 112328 6 instr_slave_r_id[7]
port 1329 nsew signal output
rlabel metal2 s 52182 359200 52238 360000 6 instr_slave_r_id[8]
port 1330 nsew signal output
rlabel metal2 s 81162 359200 81218 360000 6 instr_slave_r_id[9]
port 1331 nsew signal output
rlabel metal2 s 41234 359200 41290 360000 6 instr_slave_r_last
port 1332 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 instr_slave_r_ready
port 1333 nsew signal input
rlabel metal3 s 0 165248 800 165368 6 instr_slave_r_resp[0]
port 1334 nsew signal output
rlabel metal2 s 228638 359200 228694 360000 6 instr_slave_r_resp[1]
port 1335 nsew signal output
rlabel metal3 s 279200 58488 280000 58608 6 instr_slave_r_user[-1]
port 1336 nsew signal output
rlabel metal2 s 267278 0 267334 800 6 instr_slave_r_user[0]
port 1337 nsew signal output
rlabel metal3 s 279200 48288 280000 48408 6 instr_slave_r_valid
port 1338 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 instr_slave_w_data[0]
port 1339 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 instr_slave_w_data[10]
port 1340 nsew signal input
rlabel metal2 s 49606 359200 49662 360000 6 instr_slave_w_data[11]
port 1341 nsew signal input
rlabel metal2 s 31574 359200 31630 360000 6 instr_slave_w_data[12]
port 1342 nsew signal input
rlabel metal3 s 0 196528 800 196648 6 instr_slave_w_data[13]
port 1343 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 instr_slave_w_data[14]
port 1344 nsew signal input
rlabel metal3 s 0 325048 800 325168 6 instr_slave_w_data[15]
port 1345 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 instr_slave_w_data[16]
port 1346 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 instr_slave_w_data[17]
port 1347 nsew signal input
rlabel metal3 s 0 177488 800 177608 6 instr_slave_w_data[18]
port 1348 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 instr_slave_w_data[19]
port 1349 nsew signal input
rlabel metal3 s 279200 247528 280000 247648 6 instr_slave_w_data[1]
port 1350 nsew signal input
rlabel metal3 s 279200 233928 280000 234048 6 instr_slave_w_data[20]
port 1351 nsew signal input
rlabel metal3 s 0 223048 800 223168 6 instr_slave_w_data[21]
port 1352 nsew signal input
rlabel metal3 s 0 302608 800 302728 6 instr_slave_w_data[22]
port 1353 nsew signal input
rlabel metal2 s 104990 359200 105046 360000 6 instr_slave_w_data[23]
port 1354 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 instr_slave_w_data[24]
port 1355 nsew signal input
rlabel metal2 s 257618 359200 257674 360000 6 instr_slave_w_data[25]
port 1356 nsew signal input
rlabel metal2 s 222842 0 222898 800 6 instr_slave_w_data[26]
port 1357 nsew signal input
rlabel metal2 s 251822 0 251878 800 6 instr_slave_w_data[27]
port 1358 nsew signal input
rlabel metal2 s 220910 359200 220966 360000 6 instr_slave_w_data[28]
port 1359 nsew signal input
rlabel metal2 s 41878 359200 41934 360000 6 instr_slave_w_data[29]
port 1360 nsew signal input
rlabel metal3 s 279200 263168 280000 263288 6 instr_slave_w_data[2]
port 1361 nsew signal input
rlabel metal3 s 0 354968 800 355088 6 instr_slave_w_data[30]
port 1362 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 instr_slave_w_data[31]
port 1363 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 instr_slave_w_data[32]
port 1364 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 instr_slave_w_data[33]
port 1365 nsew signal input
rlabel metal3 s 279200 57128 280000 57248 6 instr_slave_w_data[34]
port 1366 nsew signal input
rlabel metal2 s 236366 359200 236422 360000 6 instr_slave_w_data[35]
port 1367 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 instr_slave_w_data[36]
port 1368 nsew signal input
rlabel metal2 s 76010 359200 76066 360000 6 instr_slave_w_data[37]
port 1369 nsew signal input
rlabel metal3 s 0 336608 800 336728 6 instr_slave_w_data[38]
port 1370 nsew signal input
rlabel metal3 s 279200 242768 280000 242888 6 instr_slave_w_data[39]
port 1371 nsew signal input
rlabel metal3 s 279200 106768 280000 106888 6 instr_slave_w_data[3]
port 1372 nsew signal input
rlabel metal3 s 279200 118328 280000 118448 6 instr_slave_w_data[40]
port 1373 nsew signal input
rlabel metal2 s 217690 359200 217746 360000 6 instr_slave_w_data[41]
port 1374 nsew signal input
rlabel metal3 s 0 329128 800 329248 6 instr_slave_w_data[42]
port 1375 nsew signal input
rlabel metal2 s 171966 0 172022 800 6 instr_slave_w_data[43]
port 1376 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 instr_slave_w_data[44]
port 1377 nsew signal input
rlabel metal2 s 260838 359200 260894 360000 6 instr_slave_w_data[45]
port 1378 nsew signal input
rlabel metal3 s 279200 68688 280000 68808 6 instr_slave_w_data[46]
port 1379 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 instr_slave_w_data[47]
port 1380 nsew signal input
rlabel metal2 s 96618 359200 96674 360000 6 instr_slave_w_data[48]
port 1381 nsew signal input
rlabel metal3 s 0 253648 800 253768 6 instr_slave_w_data[49]
port 1382 nsew signal input
rlabel metal2 s 193218 359200 193274 360000 6 instr_slave_w_data[4]
port 1383 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 instr_slave_w_data[50]
port 1384 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 instr_slave_w_data[51]
port 1385 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 instr_slave_w_data[52]
port 1386 nsew signal input
rlabel metal3 s 279200 47608 280000 47728 6 instr_slave_w_data[53]
port 1387 nsew signal input
rlabel metal3 s 279200 327088 280000 327208 6 instr_slave_w_data[54]
port 1388 nsew signal input
rlabel metal2 s 43166 359200 43222 360000 6 instr_slave_w_data[55]
port 1389 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 instr_slave_w_data[56]
port 1390 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 instr_slave_w_data[57]
port 1391 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 instr_slave_w_data[58]
port 1392 nsew signal input
rlabel metal3 s 279200 241408 280000 241528 6 instr_slave_w_data[59]
port 1393 nsew signal input
rlabel metal3 s 279200 43528 280000 43648 6 instr_slave_w_data[5]
port 1394 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 instr_slave_w_data[60]
port 1395 nsew signal input
rlabel metal2 s 61842 359200 61898 360000 6 instr_slave_w_data[61]
port 1396 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 instr_slave_w_data[62]
port 1397 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 instr_slave_w_data[63]
port 1398 nsew signal input
rlabel metal3 s 0 163208 800 163328 6 instr_slave_w_data[6]
port 1399 nsew signal input
rlabel metal3 s 279200 274048 280000 274168 6 instr_slave_w_data[7]
port 1400 nsew signal input
rlabel metal3 s 279200 127848 280000 127968 6 instr_slave_w_data[8]
port 1401 nsew signal input
rlabel metal2 s 262126 359200 262182 360000 6 instr_slave_w_data[9]
port 1402 nsew signal input
rlabel metal3 s 0 263848 800 263968 6 instr_slave_w_last
port 1403 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 instr_slave_w_ready
port 1404 nsew signal output
rlabel metal3 s 279200 206048 280000 206168 6 instr_slave_w_strb[0]
port 1405 nsew signal input
rlabel metal3 s 279200 97248 280000 97368 6 instr_slave_w_strb[1]
port 1406 nsew signal input
rlabel metal2 s 87602 359200 87658 360000 6 instr_slave_w_strb[2]
port 1407 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 instr_slave_w_strb[3]
port 1408 nsew signal input
rlabel metal3 s 0 229848 800 229968 6 instr_slave_w_strb[4]
port 1409 nsew signal input
rlabel metal2 s 240874 0 240930 800 6 instr_slave_w_strb[5]
port 1410 nsew signal input
rlabel metal3 s 279200 99968 280000 100088 6 instr_slave_w_strb[6]
port 1411 nsew signal input
rlabel metal2 s 126886 359200 126942 360000 6 instr_slave_w_strb[7]
port 1412 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 instr_slave_w_user[-1]
port 1413 nsew signal input
rlabel metal2 s 217046 359200 217102 360000 6 instr_slave_w_user[0]
port 1414 nsew signal input
rlabel metal3 s 279200 341368 280000 341488 6 instr_slave_w_valid
port 1415 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 irq_i[0]
port 1416 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 irq_i[10]
port 1417 nsew signal input
rlabel metal3 s 0 249568 800 249688 6 irq_i[11]
port 1418 nsew signal input
rlabel metal3 s 279200 187008 280000 187128 6 irq_i[12]
port 1419 nsew signal input
rlabel metal3 s 279200 232568 280000 232688 6 irq_i[13]
port 1420 nsew signal input
rlabel metal3 s 0 207408 800 207528 6 irq_i[14]
port 1421 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 irq_i[15]
port 1422 nsew signal input
rlabel metal2 s 204166 359200 204222 360000 6 irq_i[16]
port 1423 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 irq_i[17]
port 1424 nsew signal input
rlabel metal2 s 251178 359200 251234 360000 6 irq_i[18]
port 1425 nsew signal input
rlabel metal3 s 0 327088 800 327208 6 irq_i[19]
port 1426 nsew signal input
rlabel metal3 s 0 202648 800 202768 6 irq_i[1]
port 1427 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 irq_i[20]
port 1428 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 irq_i[21]
port 1429 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 irq_i[22]
port 1430 nsew signal input
rlabel metal3 s 279200 150968 280000 151088 6 irq_i[23]
port 1431 nsew signal input
rlabel metal3 s 279200 250248 280000 250368 6 irq_i[24]
port 1432 nsew signal input
rlabel metal3 s 0 248208 800 248328 6 irq_i[25]
port 1433 nsew signal input
rlabel metal2 s 271786 359200 271842 360000 6 irq_i[26]
port 1434 nsew signal input
rlabel metal2 s 275006 0 275062 800 6 irq_i[27]
port 1435 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 irq_i[28]
port 1436 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 irq_i[29]
port 1437 nsew signal input
rlabel metal3 s 279200 14968 280000 15088 6 irq_i[2]
port 1438 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 irq_i[30]
port 1439 nsew signal input
rlabel metal3 s 279200 33328 280000 33448 6 irq_i[31]
port 1440 nsew signal input
rlabel metal2 s 162306 359200 162362 360000 6 irq_i[3]
port 1441 nsew signal input
rlabel metal3 s 279200 248888 280000 249008 6 irq_i[4]
port 1442 nsew signal input
rlabel metal2 s 178406 359200 178462 360000 6 irq_i[5]
port 1443 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 irq_i[6]
port 1444 nsew signal input
rlabel metal3 s 0 203328 800 203448 6 irq_i[7]
port 1445 nsew signal input
rlabel metal3 s 0 254328 800 254448 6 irq_i[8]
port 1446 nsew signal input
rlabel metal2 s 264058 0 264114 800 6 irq_i[9]
port 1447 nsew signal input
rlabel metal3 s 0 242088 800 242208 6 mba_data_mem_addr0_o[0]
port 1448 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 mba_data_mem_addr0_o[10]
port 1449 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 mba_data_mem_addr0_o[11]
port 1450 nsew signal output
rlabel metal3 s 279200 148928 280000 149048 6 mba_data_mem_addr0_o[12]
port 1451 nsew signal output
rlabel metal2 s 166814 359200 166870 360000 6 mba_data_mem_addr0_o[13]
port 1452 nsew signal output
rlabel metal3 s 279200 319608 280000 319728 6 mba_data_mem_addr0_o[14]
port 1453 nsew signal output
rlabel metal3 s 279200 277448 280000 277568 6 mba_data_mem_addr0_o[15]
port 1454 nsew signal output
rlabel metal2 s 228638 0 228694 800 6 mba_data_mem_addr0_o[16]
port 1455 nsew signal output
rlabel metal3 s 279200 61208 280000 61328 6 mba_data_mem_addr0_o[17]
port 1456 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 mba_data_mem_addr0_o[18]
port 1457 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 mba_data_mem_addr0_o[19]
port 1458 nsew signal output
rlabel metal2 s 256330 0 256386 800 6 mba_data_mem_addr0_o[1]
port 1459 nsew signal output
rlabel metal3 s 279200 78208 280000 78328 6 mba_data_mem_addr0_o[20]
port 1460 nsew signal output
rlabel metal3 s 0 144168 800 144288 6 mba_data_mem_addr0_o[21]
port 1461 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 mba_data_mem_addr0_o[22]
port 1462 nsew signal output
rlabel metal2 s 171966 359200 172022 360000 6 mba_data_mem_addr0_o[23]
port 1463 nsew signal output
rlabel metal2 s 233790 0 233846 800 6 mba_data_mem_addr0_o[24]
port 1464 nsew signal output
rlabel metal3 s 279200 243448 280000 243568 6 mba_data_mem_addr0_o[25]
port 1465 nsew signal output
rlabel metal3 s 279200 168648 280000 168768 6 mba_data_mem_addr0_o[26]
port 1466 nsew signal output
rlabel metal3 s 279200 299208 280000 299328 6 mba_data_mem_addr0_o[27]
port 1467 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 mba_data_mem_addr0_o[28]
port 1468 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 mba_data_mem_addr0_o[29]
port 1469 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 mba_data_mem_addr0_o[2]
port 1470 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 mba_data_mem_addr0_o[30]
port 1471 nsew signal output
rlabel metal3 s 0 349528 800 349648 6 mba_data_mem_addr0_o[31]
port 1472 nsew signal output
rlabel metal3 s 279200 98608 280000 98728 6 mba_data_mem_addr0_o[3]
port 1473 nsew signal output
rlabel metal2 s 33506 359200 33562 360000 6 mba_data_mem_addr0_o[4]
port 1474 nsew signal output
rlabel metal2 s 18 0 74 800 6 mba_data_mem_addr0_o[5]
port 1475 nsew signal output
rlabel metal3 s 279200 182928 280000 183048 6 mba_data_mem_addr0_o[6]
port 1476 nsew signal output
rlabel metal2 s 213182 359200 213238 360000 6 mba_data_mem_addr0_o[7]
port 1477 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 mba_data_mem_addr0_o[8]
port 1478 nsew signal output
rlabel metal3 s 279200 9528 280000 9648 6 mba_data_mem_addr0_o[9]
port 1479 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 mba_data_mem_addr1_o[0]
port 1480 nsew signal output
rlabel metal3 s 0 291048 800 291168 6 mba_data_mem_addr1_o[10]
port 1481 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 mba_data_mem_addr1_o[11]
port 1482 nsew signal output
rlabel metal3 s 279200 105408 280000 105528 6 mba_data_mem_addr1_o[12]
port 1483 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 mba_data_mem_addr1_o[13]
port 1484 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 mba_data_mem_addr1_o[14]
port 1485 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 mba_data_mem_addr1_o[15]
port 1486 nsew signal output
rlabel metal3 s 279200 70048 280000 70168 6 mba_data_mem_addr1_o[16]
port 1487 nsew signal output
rlabel metal3 s 279200 313488 280000 313608 6 mba_data_mem_addr1_o[17]
port 1488 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 mba_data_mem_addr1_o[18]
port 1489 nsew signal output
rlabel metal3 s 0 301248 800 301368 6 mba_data_mem_addr1_o[19]
port 1490 nsew signal output
rlabel metal3 s 0 161848 800 161968 6 mba_data_mem_addr1_o[1]
port 1491 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 mba_data_mem_addr1_o[20]
port 1492 nsew signal output
rlabel metal2 s 234434 0 234490 800 6 mba_data_mem_addr1_o[21]
port 1493 nsew signal output
rlabel metal2 s 37370 359200 37426 360000 6 mba_data_mem_addr1_o[22]
port 1494 nsew signal output
rlabel metal3 s 279200 222368 280000 222488 6 mba_data_mem_addr1_o[23]
port 1495 nsew signal output
rlabel metal3 s 0 320968 800 321088 6 mba_data_mem_addr1_o[24]
port 1496 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 mba_data_mem_addr1_o[25]
port 1497 nsew signal output
rlabel metal2 s 218334 359200 218390 360000 6 mba_data_mem_addr1_o[26]
port 1498 nsew signal output
rlabel metal3 s 279200 40808 280000 40928 6 mba_data_mem_addr1_o[27]
port 1499 nsew signal output
rlabel metal2 s 28354 359200 28410 360000 6 mba_data_mem_addr1_o[28]
port 1500 nsew signal output
rlabel metal2 s 226706 359200 226762 360000 6 mba_data_mem_addr1_o[29]
port 1501 nsew signal output
rlabel metal3 s 0 250928 800 251048 6 mba_data_mem_addr1_o[2]
port 1502 nsew signal output
rlabel metal3 s 0 306008 800 306128 6 mba_data_mem_addr1_o[30]
port 1503 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 mba_data_mem_addr1_o[31]
port 1504 nsew signal output
rlabel metal2 s 148782 359200 148838 360000 6 mba_data_mem_addr1_o[3]
port 1505 nsew signal output
rlabel metal3 s 279200 35368 280000 35488 6 mba_data_mem_addr1_o[4]
port 1506 nsew signal output
rlabel metal2 s 251822 359200 251878 360000 6 mba_data_mem_addr1_o[5]
port 1507 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 mba_data_mem_addr1_o[6]
port 1508 nsew signal output
rlabel metal3 s 0 230528 800 230648 6 mba_data_mem_addr1_o[7]
port 1509 nsew signal output
rlabel metal2 s 247958 0 248014 800 6 mba_data_mem_addr1_o[8]
port 1510 nsew signal output
rlabel metal2 s 220266 0 220322 800 6 mba_data_mem_addr1_o[9]
port 1511 nsew signal output
rlabel metal2 s 79230 359200 79286 360000 6 mba_data_mem_csb0_o
port 1512 nsew signal output
rlabel metal3 s 279200 324368 280000 324488 6 mba_data_mem_csb1_o
port 1513 nsew signal output
rlabel metal3 s 279200 176128 280000 176248 6 mba_data_mem_din0_o[0]
port 1514 nsew signal output
rlabel metal2 s 242162 359200 242218 360000 6 mba_data_mem_din0_o[10]
port 1515 nsew signal output
rlabel metal2 s 271142 0 271198 800 6 mba_data_mem_din0_o[11]
port 1516 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 mba_data_mem_din0_o[12]
port 1517 nsew signal output
rlabel metal3 s 0 265208 800 265328 6 mba_data_mem_din0_o[13]
port 1518 nsew signal output
rlabel metal2 s 141054 359200 141110 360000 6 mba_data_mem_din0_o[14]
port 1519 nsew signal output
rlabel metal3 s 279200 291728 280000 291848 6 mba_data_mem_din0_o[15]
port 1520 nsew signal output
rlabel metal3 s 279200 354968 280000 355088 6 mba_data_mem_din0_o[16]
port 1521 nsew signal output
rlabel metal3 s 279200 67328 280000 67448 6 mba_data_mem_din0_o[17]
port 1522 nsew signal output
rlabel metal3 s 279200 253648 280000 253768 6 mba_data_mem_din0_o[18]
port 1523 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 mba_data_mem_din0_o[19]
port 1524 nsew signal output
rlabel metal3 s 0 273368 800 273488 6 mba_data_mem_din0_o[1]
port 1525 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 mba_data_mem_din0_o[20]
port 1526 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 mba_data_mem_din0_o[21]
port 1527 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 mba_data_mem_din0_o[22]
port 1528 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 mba_data_mem_din0_o[23]
port 1529 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 mba_data_mem_din0_o[24]
port 1530 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 mba_data_mem_din0_o[25]
port 1531 nsew signal output
rlabel metal3 s 279200 201288 280000 201408 6 mba_data_mem_din0_o[26]
port 1532 nsew signal output
rlabel metal2 s 117226 359200 117282 360000 6 mba_data_mem_din0_o[27]
port 1533 nsew signal output
rlabel metal3 s 279200 312808 280000 312928 6 mba_data_mem_din0_o[28]
port 1534 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 mba_data_mem_din0_o[29]
port 1535 nsew signal output
rlabel metal3 s 279200 280168 280000 280288 6 mba_data_mem_din0_o[2]
port 1536 nsew signal output
rlabel metal3 s 279200 2728 280000 2848 6 mba_data_mem_din0_o[30]
port 1537 nsew signal output
rlabel metal2 s 47674 359200 47730 360000 6 mba_data_mem_din0_o[31]
port 1538 nsew signal output
rlabel metal2 s 260838 0 260894 800 6 mba_data_mem_din0_o[3]
port 1539 nsew signal output
rlabel metal2 s 278870 359200 278926 360000 6 mba_data_mem_din0_o[4]
port 1540 nsew signal output
rlabel metal2 s 100482 359200 100538 360000 6 mba_data_mem_din0_o[5]
port 1541 nsew signal output
rlabel metal2 s 56690 359200 56746 360000 6 mba_data_mem_din0_o[6]
port 1542 nsew signal output
rlabel metal3 s 0 316888 800 317008 6 mba_data_mem_din0_o[7]
port 1543 nsew signal output
rlabel metal2 s 108210 359200 108266 360000 6 mba_data_mem_din0_o[8]
port 1544 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 mba_data_mem_din0_o[9]
port 1545 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 mba_data_mem_dout0_i[0]
port 1546 nsew signal input
rlabel metal3 s 279200 153688 280000 153808 6 mba_data_mem_dout0_i[10]
port 1547 nsew signal input
rlabel metal3 s 279200 259088 280000 259208 6 mba_data_mem_dout0_i[11]
port 1548 nsew signal input
rlabel metal2 s 275650 359200 275706 360000 6 mba_data_mem_dout0_i[12]
port 1549 nsew signal input
rlabel metal3 s 0 266568 800 266688 6 mba_data_mem_dout0_i[13]
port 1550 nsew signal input
rlabel metal3 s 279200 27888 280000 28008 6 mba_data_mem_dout0_i[14]
port 1551 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 mba_data_mem_dout0_i[15]
port 1552 nsew signal input
rlabel metal2 s 240230 359200 240286 360000 6 mba_data_mem_dout0_i[16]
port 1553 nsew signal input
rlabel metal2 s 85670 359200 85726 360000 6 mba_data_mem_dout0_i[17]
port 1554 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 mba_data_mem_dout0_i[18]
port 1555 nsew signal input
rlabel metal3 s 279200 87728 280000 87848 6 mba_data_mem_dout0_i[19]
port 1556 nsew signal input
rlabel metal2 s 151358 359200 151414 360000 6 mba_data_mem_dout0_i[1]
port 1557 nsew signal input
rlabel metal3 s 279200 72088 280000 72208 6 mba_data_mem_dout0_i[20]
port 1558 nsew signal input
rlabel metal3 s 279200 143488 280000 143608 6 mba_data_mem_dout0_i[21]
port 1559 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 mba_data_mem_dout0_i[22]
port 1560 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 mba_data_mem_dout0_i[23]
port 1561 nsew signal input
rlabel metal3 s 279200 95888 280000 96008 6 mba_data_mem_dout0_i[24]
port 1562 nsew signal input
rlabel metal3 s 279200 237328 280000 237448 6 mba_data_mem_dout0_i[25]
port 1563 nsew signal input
rlabel metal2 s 199658 359200 199714 360000 6 mba_data_mem_dout0_i[26]
port 1564 nsew signal input
rlabel metal3 s 0 300568 800 300688 6 mba_data_mem_dout0_i[27]
port 1565 nsew signal input
rlabel metal3 s 0 284928 800 285048 6 mba_data_mem_dout0_i[28]
port 1566 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 mba_data_mem_dout0_i[29]
port 1567 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 mba_data_mem_dout0_i[2]
port 1568 nsew signal input
rlabel metal2 s 166170 359200 166226 360000 6 mba_data_mem_dout0_i[30]
port 1569 nsew signal input
rlabel metal3 s 279200 131248 280000 131368 6 mba_data_mem_dout0_i[31]
port 1570 nsew signal input
rlabel metal3 s 0 206048 800 206168 6 mba_data_mem_dout0_i[3]
port 1571 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 mba_data_mem_dout0_i[4]
port 1572 nsew signal input
rlabel metal2 s 215114 359200 215170 360000 6 mba_data_mem_dout0_i[5]
port 1573 nsew signal input
rlabel metal2 s 27710 359200 27766 360000 6 mba_data_mem_dout0_i[6]
port 1574 nsew signal input
rlabel metal2 s 5170 359200 5226 360000 6 mba_data_mem_dout0_i[7]
port 1575 nsew signal input
rlabel metal2 s 74722 359200 74778 360000 6 mba_data_mem_dout0_i[8]
port 1576 nsew signal input
rlabel metal2 s 94042 359200 94098 360000 6 mba_data_mem_dout0_i[9]
port 1577 nsew signal input
rlabel metal2 s 98550 359200 98606 360000 6 mba_data_mem_web0_o
port 1578 nsew signal output
rlabel metal2 s 224774 0 224830 800 6 mba_data_mem_wmask0_o[0]
port 1579 nsew signal output
rlabel metal3 s 0 332528 800 332648 6 mba_data_mem_wmask0_o[1]
port 1580 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 mba_data_mem_wmask0_o[2]
port 1581 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 mba_data_mem_wmask0_o[3]
port 1582 nsew signal output
rlabel metal3 s 279200 56448 280000 56568 6 mba_instr_mem_addr0_o[0]
port 1583 nsew signal output
rlabel metal2 s 226062 0 226118 800 6 mba_instr_mem_addr0_o[10]
port 1584 nsew signal output
rlabel metal3 s 279200 178848 280000 178968 6 mba_instr_mem_addr0_o[11]
port 1585 nsew signal output
rlabel metal2 s 19982 359200 20038 360000 6 mba_instr_mem_addr0_o[12]
port 1586 nsew signal output
rlabel metal3 s 279200 214208 280000 214328 6 mba_instr_mem_addr0_o[13]
port 1587 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 mba_instr_mem_addr0_o[14]
port 1588 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 mba_instr_mem_addr0_o[15]
port 1589 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 mba_instr_mem_addr0_o[16]
port 1590 nsew signal output
rlabel metal2 s 188066 0 188122 800 6 mba_instr_mem_addr0_o[17]
port 1591 nsew signal output
rlabel metal3 s 0 341368 800 341488 6 mba_instr_mem_addr0_o[18]
port 1592 nsew signal output
rlabel metal3 s 279200 61888 280000 62008 6 mba_instr_mem_addr0_o[19]
port 1593 nsew signal output
rlabel metal2 s 161018 0 161074 800 6 mba_instr_mem_addr0_o[1]
port 1594 nsew signal output
rlabel metal3 s 279200 38768 280000 38888 6 mba_instr_mem_addr0_o[20]
port 1595 nsew signal output
rlabel metal2 s 277582 359200 277638 360000 6 mba_instr_mem_addr0_o[21]
port 1596 nsew signal output
rlabel metal2 s 203522 359200 203578 360000 6 mba_instr_mem_addr0_o[22]
port 1597 nsew signal output
rlabel metal3 s 279200 44208 280000 44328 6 mba_instr_mem_addr0_o[23]
port 1598 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 mba_instr_mem_addr0_o[24]
port 1599 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 mba_instr_mem_addr0_o[25]
port 1600 nsew signal output
rlabel metal2 s 225418 359200 225474 360000 6 mba_instr_mem_addr0_o[26]
port 1601 nsew signal output
rlabel metal3 s 0 303288 800 303408 6 mba_instr_mem_addr0_o[27]
port 1602 nsew signal output
rlabel metal2 s 278226 359200 278282 360000 6 mba_instr_mem_addr0_o[28]
port 1603 nsew signal output
rlabel metal3 s 279200 34688 280000 34808 6 mba_instr_mem_addr0_o[29]
port 1604 nsew signal output
rlabel metal2 s 38014 359200 38070 360000 6 mba_instr_mem_addr0_o[2]
port 1605 nsew signal output
rlabel metal3 s 279200 178168 280000 178288 6 mba_instr_mem_addr0_o[30]
port 1606 nsew signal output
rlabel metal3 s 0 280168 800 280288 6 mba_instr_mem_addr0_o[31]
port 1607 nsew signal output
rlabel metal3 s 279200 101328 280000 101448 6 mba_instr_mem_addr0_o[3]
port 1608 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 mba_instr_mem_addr0_o[4]
port 1609 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 mba_instr_mem_addr0_o[5]
port 1610 nsew signal output
rlabel metal3 s 279200 342048 280000 342168 6 mba_instr_mem_addr0_o[6]
port 1611 nsew signal output
rlabel metal2 s 226706 0 226762 800 6 mba_instr_mem_addr0_o[7]
port 1612 nsew signal output
rlabel metal2 s 238942 359200 238998 360000 6 mba_instr_mem_addr0_o[8]
port 1613 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 mba_instr_mem_addr0_o[9]
port 1614 nsew signal output
rlabel metal3 s 279200 104728 280000 104848 6 mba_instr_mem_addr1_o[0]
port 1615 nsew signal output
rlabel metal3 s 0 180208 800 180328 6 mba_instr_mem_addr1_o[10]
port 1616 nsew signal output
rlabel metal2 s 55402 359200 55458 360000 6 mba_instr_mem_addr1_o[11]
port 1617 nsew signal output
rlabel metal2 s 204810 359200 204866 360000 6 mba_instr_mem_addr1_o[12]
port 1618 nsew signal output
rlabel metal3 s 0 171368 800 171488 6 mba_instr_mem_addr1_o[13]
port 1619 nsew signal output
rlabel metal3 s 0 210128 800 210248 6 mba_instr_mem_addr1_o[14]
port 1620 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 mba_instr_mem_addr1_o[15]
port 1621 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 mba_instr_mem_addr1_o[16]
port 1622 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 mba_instr_mem_addr1_o[17]
port 1623 nsew signal output
rlabel metal3 s 0 355648 800 355768 6 mba_instr_mem_addr1_o[18]
port 1624 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 mba_instr_mem_addr1_o[19]
port 1625 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 mba_instr_mem_addr1_o[1]
port 1626 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 mba_instr_mem_addr1_o[20]
port 1627 nsew signal output
rlabel metal2 s 215758 0 215814 800 6 mba_instr_mem_addr1_o[21]
port 1628 nsew signal output
rlabel metal2 s 235722 359200 235778 360000 6 mba_instr_mem_addr1_o[22]
port 1629 nsew signal output
rlabel metal2 s 259550 359200 259606 360000 6 mba_instr_mem_addr1_o[23]
port 1630 nsew signal output
rlabel metal2 s 244094 0 244150 800 6 mba_instr_mem_addr1_o[24]
port 1631 nsew signal output
rlabel metal3 s 279200 348848 280000 348968 6 mba_instr_mem_addr1_o[25]
port 1632 nsew signal output
rlabel metal3 s 279200 231888 280000 232008 6 mba_instr_mem_addr1_o[26]
port 1633 nsew signal output
rlabel metal3 s 279200 91128 280000 91248 6 mba_instr_mem_addr1_o[27]
port 1634 nsew signal output
rlabel metal2 s 12254 359200 12310 360000 6 mba_instr_mem_addr1_o[28]
port 1635 nsew signal output
rlabel metal2 s 121090 359200 121146 360000 6 mba_instr_mem_addr1_o[29]
port 1636 nsew signal output
rlabel metal2 s 214470 0 214526 800 6 mba_instr_mem_addr1_o[2]
port 1637 nsew signal output
rlabel metal3 s 279200 25168 280000 25288 6 mba_instr_mem_addr1_o[30]
port 1638 nsew signal output
rlabel metal3 s 279200 190408 280000 190528 6 mba_instr_mem_addr1_o[31]
port 1639 nsew signal output
rlabel metal3 s 0 178168 800 178288 6 mba_instr_mem_addr1_o[3]
port 1640 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 mba_instr_mem_addr1_o[4]
port 1641 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 mba_instr_mem_addr1_o[5]
port 1642 nsew signal output
rlabel metal3 s 0 272008 800 272128 6 mba_instr_mem_addr1_o[6]
port 1643 nsew signal output
rlabel metal3 s 279200 323008 280000 323128 6 mba_instr_mem_addr1_o[7]
port 1644 nsew signal output
rlabel metal2 s 179050 359200 179106 360000 6 mba_instr_mem_addr1_o[8]
port 1645 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 mba_instr_mem_addr1_o[9]
port 1646 nsew signal output
rlabel metal2 s 91466 359200 91522 360000 6 mba_instr_mem_csb0_o
port 1647 nsew signal output
rlabel metal3 s 279200 255008 280000 255128 6 mba_instr_mem_csb1_o
port 1648 nsew signal output
rlabel metal3 s 279200 5448 280000 5568 6 mba_instr_mem_din0_o[0]
port 1649 nsew signal output
rlabel metal2 s 88890 359200 88946 360000 6 mba_instr_mem_din0_o[10]
port 1650 nsew signal output
rlabel metal2 s 274362 0 274418 800 6 mba_instr_mem_din0_o[11]
port 1651 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 mba_instr_mem_din0_o[12]
port 1652 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 mba_instr_mem_din0_o[13]
port 1653 nsew signal output
rlabel metal3 s 279200 86368 280000 86488 6 mba_instr_mem_din0_o[14]
port 1654 nsew signal output
rlabel metal3 s 279200 188368 280000 188488 6 mba_instr_mem_din0_o[15]
port 1655 nsew signal output
rlabel metal3 s 0 294448 800 294568 6 mba_instr_mem_din0_o[16]
port 1656 nsew signal output
rlabel metal2 s 229282 359200 229338 360000 6 mba_instr_mem_din0_o[17]
port 1657 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 mba_instr_mem_din0_o[18]
port 1658 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 mba_instr_mem_din0_o[19]
port 1659 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 mba_instr_mem_din0_o[1]
port 1660 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 mba_instr_mem_din0_o[20]
port 1661 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 mba_instr_mem_din0_o[21]
port 1662 nsew signal output
rlabel metal3 s 279200 273368 280000 273488 6 mba_instr_mem_din0_o[22]
port 1663 nsew signal output
rlabel metal2 s 203522 0 203578 800 6 mba_instr_mem_din0_o[23]
port 1664 nsew signal output
rlabel metal2 s 86314 359200 86370 360000 6 mba_instr_mem_din0_o[24]
port 1665 nsew signal output
rlabel metal2 s 172610 359200 172666 360000 6 mba_instr_mem_din0_o[25]
port 1666 nsew signal output
rlabel metal3 s 0 222368 800 222488 6 mba_instr_mem_din0_o[26]
port 1667 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 mba_instr_mem_din0_o[27]
port 1668 nsew signal output
rlabel metal3 s 279200 296488 280000 296608 6 mba_instr_mem_din0_o[28]
port 1669 nsew signal output
rlabel metal2 s 189354 359200 189410 360000 6 mba_instr_mem_din0_o[29]
port 1670 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 mba_instr_mem_din0_o[2]
port 1671 nsew signal output
rlabel metal3 s 279200 357008 280000 357128 6 mba_instr_mem_din0_o[30]
port 1672 nsew signal output
rlabel metal3 s 279200 189728 280000 189848 6 mba_instr_mem_din0_o[31]
port 1673 nsew signal output
rlabel metal2 s 240230 0 240286 800 6 mba_instr_mem_din0_o[3]
port 1674 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 mba_instr_mem_din0_o[4]
port 1675 nsew signal output
rlabel metal3 s 0 312128 800 312248 6 mba_instr_mem_din0_o[5]
port 1676 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 mba_instr_mem_din0_o[6]
port 1677 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 mba_instr_mem_din0_o[7]
port 1678 nsew signal output
rlabel metal3 s 279200 688 280000 808 6 mba_instr_mem_din0_o[8]
port 1679 nsew signal output
rlabel metal3 s 279200 171368 280000 171488 6 mba_instr_mem_din0_o[9]
port 1680 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 mba_instr_mem_dout0_i[0]
port 1681 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 mba_instr_mem_dout0_i[10]
port 1682 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 mba_instr_mem_dout0_i[11]
port 1683 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 mba_instr_mem_dout0_i[12]
port 1684 nsew signal input
rlabel metal3 s 279200 215568 280000 215688 6 mba_instr_mem_dout0_i[13]
port 1685 nsew signal input
rlabel metal2 s 159086 359200 159142 360000 6 mba_instr_mem_dout0_i[14]
port 1686 nsew signal input
rlabel metal2 s 264058 359200 264114 360000 6 mba_instr_mem_dout0_i[15]
port 1687 nsew signal input
rlabel metal3 s 279200 77528 280000 77648 6 mba_instr_mem_dout0_i[16]
port 1688 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 mba_instr_mem_dout0_i[17]
port 1689 nsew signal input
rlabel metal3 s 279200 258408 280000 258528 6 mba_instr_mem_dout0_i[18]
port 1690 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 mba_instr_mem_dout0_i[19]
port 1691 nsew signal input
rlabel metal2 s 262770 359200 262826 360000 6 mba_instr_mem_dout0_i[1]
port 1692 nsew signal input
rlabel metal2 s 155866 359200 155922 360000 6 mba_instr_mem_dout0_i[20]
port 1693 nsew signal input
rlabel metal3 s 279200 95208 280000 95328 6 mba_instr_mem_dout0_i[21]
port 1694 nsew signal input
rlabel metal2 s 148138 359200 148194 360000 6 mba_instr_mem_dout0_i[22]
port 1695 nsew signal input
rlabel metal2 s 223486 0 223542 800 6 mba_instr_mem_dout0_i[23]
port 1696 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 mba_instr_mem_dout0_i[24]
port 1697 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 mba_instr_mem_dout0_i[25]
port 1698 nsew signal input
rlabel metal2 s 662 0 718 800 6 mba_instr_mem_dout0_i[26]
port 1699 nsew signal input
rlabel metal2 s 258906 0 258962 800 6 mba_instr_mem_dout0_i[27]
port 1700 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 mba_instr_mem_dout0_i[28]
port 1701 nsew signal input
rlabel metal3 s 0 235288 800 235408 6 mba_instr_mem_dout0_i[29]
port 1702 nsew signal input
rlabel metal2 s 16118 359200 16174 360000 6 mba_instr_mem_dout0_i[2]
port 1703 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 mba_instr_mem_dout0_i[30]
port 1704 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 mba_instr_mem_dout0_i[31]
port 1705 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 mba_instr_mem_dout0_i[3]
port 1706 nsew signal input
rlabel metal2 s 101126 359200 101182 360000 6 mba_instr_mem_dout0_i[4]
port 1707 nsew signal input
rlabel metal2 s 30930 359200 30986 360000 6 mba_instr_mem_dout0_i[5]
port 1708 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 mba_instr_mem_dout0_i[6]
port 1709 nsew signal input
rlabel metal2 s 161662 359200 161718 360000 6 mba_instr_mem_dout0_i[7]
port 1710 nsew signal input
rlabel metal3 s 279200 137368 280000 137488 6 mba_instr_mem_dout0_i[8]
port 1711 nsew signal input
rlabel metal3 s 0 184968 800 185088 6 mba_instr_mem_dout0_i[9]
port 1712 nsew signal input
rlabel metal3 s 279200 301248 280000 301368 6 mba_instr_mem_web0_o
port 1713 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 mba_instr_mem_wmask0_o[0]
port 1714 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 mba_instr_mem_wmask0_o[1]
port 1715 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 mba_instr_mem_wmask0_o[2]
port 1716 nsew signal output
rlabel metal3 s 279200 285608 280000 285728 6 mba_instr_mem_wmask0_o[3]
port 1717 nsew signal output
rlabel metal2 s 192574 0 192630 800 6 rst_n
port 1718 nsew signal input
rlabel metal2 s 162950 359200 163006 360000 6 tck_i
port 1719 nsew signal input
rlabel metal2 s 160374 359200 160430 360000 6 tdi_i
port 1720 nsew signal input
rlabel metal3 s 0 292408 800 292528 6 tdo_o
port 1721 nsew signal output
rlabel metal3 s 0 354288 800 354408 6 testmode_i
port 1722 nsew signal input
rlabel metal2 s 227350 0 227406 800 6 tms_i
port 1723 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 trstn_i
port 1724 nsew signal input
rlabel metal3 s 0 267248 800 267368 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 357456 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal4 s 34928 2128 35248 357456 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal4 s 65648 2128 65968 357456 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal4 s 96368 2128 96688 357456 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal4 s 127088 2128 127408 357456 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal4 s 157808 2128 158128 357456 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal4 s 188528 2128 188848 357456 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal4 s 219248 2128 219568 357456 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal4 s 249968 2128 250288 357456 6 vccd1
port 1725 nsew signal bidirectional
rlabel metal3 s 279200 195168 280000 195288 6 vssd1
port 1726 nsew signal bidirectional
rlabel metal4 s 19568 2128 19888 357456 6 vssd1
port 1726 nsew signal bidirectional
rlabel metal4 s 50288 2128 50608 357456 6 vssd1
port 1726 nsew signal bidirectional
rlabel metal4 s 81008 2128 81328 357456 6 vssd1
port 1726 nsew signal bidirectional
rlabel metal4 s 111728 2128 112048 357456 6 vssd1
port 1726 nsew signal bidirectional
rlabel metal4 s 142448 2128 142768 357456 6 vssd1
port 1726 nsew signal bidirectional
rlabel metal4 s 173168 2128 173488 357456 6 vssd1
port 1726 nsew signal bidirectional
rlabel metal4 s 203888 2128 204208 357456 6 vssd1
port 1726 nsew signal bidirectional
rlabel metal4 s 234608 2128 234928 357456 6 vssd1
port 1726 nsew signal bidirectional
rlabel metal4 s 265328 2128 265648 357456 6 vssd1
port 1726 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 280000 360000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 106957278
string GDS_FILE /home/mbaykenar/Desktop/workspace/mpw7_yonga_soc/openlane/mba_core_region/runs/22_08_03_22_53/results/signoff/mba_core_region.magic.gds
string GDS_START 1728280
<< end >>

